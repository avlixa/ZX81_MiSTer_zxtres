-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Alastair M. Robinson for the ZPUFlex project.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.zpupkg.all;

entity CtrlROM_ROM is
generic
	(
		maxAddrBitBRAM : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_zpu : in ZPU_ToROM;
	to_zpu : out ZPU_FromROM
);
end CtrlROM_ROM;

architecture arch of CtrlROM_ROM is

type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"0b0b0b0b",
     1 => x"8c0b0b0b",
     2 => x"0b81e004",
     3 => x"0b0b0b0b",
     4 => x"8c04ff0d",
     5 => x"80040400",
     6 => x"00000016",
     7 => x"00000000",
     8 => x"0b0b80dd",
     9 => x"cc080b0b",
    10 => x"80ddd008",
    11 => x"0b0b80dd",
    12 => x"d4080b0b",
    13 => x"0b0b9808",
    14 => x"2d0b0b80",
    15 => x"ddd40c0b",
    16 => x"0b80ddd0",
    17 => x"0c0b0b80",
    18 => x"ddcc0c04",
    19 => x"00000000",
    20 => x"00000000",
    21 => x"00000000",
    22 => x"00000000",
    23 => x"00000000",
    24 => x"71fd0608",
    25 => x"72830609",
    26 => x"81058205",
    27 => x"832b2a83",
    28 => x"ffff0652",
    29 => x"0471fc06",
    30 => x"08728306",
    31 => x"09810583",
    32 => x"05101010",
    33 => x"2a81ff06",
    34 => x"520471fd",
    35 => x"060883ff",
    36 => x"ff738306",
    37 => x"09810582",
    38 => x"05832b2b",
    39 => x"09067383",
    40 => x"ffff0673",
    41 => x"83060981",
    42 => x"05820583",
    43 => x"2b0b2b07",
    44 => x"72fc060c",
    45 => x"51510471",
    46 => x"fc06080b",
    47 => x"0b80c6a8",
    48 => x"73830610",
    49 => x"10050806",
    50 => x"7381ff06",
    51 => x"73830609",
    52 => x"81058305",
    53 => x"1010102b",
    54 => x"0772fc06",
    55 => x"0c515104",
    56 => x"80ddcc70",
    57 => x"80ea9027",
    58 => x"8b388071",
    59 => x"70840553",
    60 => x"0c81e304",
    61 => x"8c519089",
    62 => x"0402fc05",
    63 => x"0df88051",
    64 => x"8f0b80dd",
    65 => x"dc0c9f0b",
    66 => x"80dde00c",
    67 => x"a0717081",
    68 => x"05533480",
    69 => x"dde008ff",
    70 => x"0580dde0",
    71 => x"0c80dde0",
    72 => x"088025e8",
    73 => x"3880dddc",
    74 => x"08ff0580",
    75 => x"dddc0c80",
    76 => x"dddc0880",
    77 => x"25d03880",
    78 => x"0b80dde0",
    79 => x"0c800b80",
    80 => x"dddc0c02",
    81 => x"84050d04",
    82 => x"02f0050d",
    83 => x"f88053f8",
    84 => x"a05483bf",
    85 => x"52737081",
    86 => x"05553351",
    87 => x"70737081",
    88 => x"055534ff",
    89 => x"12527180",
    90 => x"25eb38fb",
    91 => x"c0539f52",
    92 => x"a0737081",
    93 => x"055534ff",
    94 => x"12527180",
    95 => x"25f23802",
    96 => x"90050d04",
    97 => x"02f4050d",
    98 => x"74538e0b",
    99 => x"80dddc08",
   100 => x"25913882",
   101 => x"c82d80dd",
   102 => x"dc08ff05",
   103 => x"80dddc0c",
   104 => x"838a0480",
   105 => x"dddc0880",
   106 => x"dde00853",
   107 => x"51728a2e",
   108 => x"098106be",
   109 => x"38715171",
   110 => x"9f24a438",
   111 => x"80dddc08",
   112 => x"a02911f8",
   113 => x"80115151",
   114 => x"a0713480",
   115 => x"dde00881",
   116 => x"0580dde0",
   117 => x"0c80dde0",
   118 => x"08519f71",
   119 => x"25de3880",
   120 => x"0b80dde0",
   121 => x"0c80dddc",
   122 => x"08810580",
   123 => x"dddc0c84",
   124 => x"880470a0",
   125 => x"2912f880",
   126 => x"11515172",
   127 => x"713480dd",
   128 => x"e0088105",
   129 => x"80dde00c",
   130 => x"80dde008",
   131 => x"a02e0981",
   132 => x"06913880",
   133 => x"0b80dde0",
   134 => x"0c80dddc",
   135 => x"08810580",
   136 => x"dddc0c02",
   137 => x"8c050d04",
   138 => x"02e8050d",
   139 => x"77795656",
   140 => x"880bfc16",
   141 => x"77712c8f",
   142 => x"06545254",
   143 => x"80537272",
   144 => x"25953871",
   145 => x"53fbe014",
   146 => x"51877134",
   147 => x"8114ff14",
   148 => x"545472f1",
   149 => x"387153f9",
   150 => x"1576712c",
   151 => x"87065351",
   152 => x"71802e8b",
   153 => x"38fbe014",
   154 => x"51717134",
   155 => x"81145472",
   156 => x"8e249538",
   157 => x"8f733153",
   158 => x"fbe01451",
   159 => x"a0713481",
   160 => x"14ff1454",
   161 => x"5472f138",
   162 => x"0298050d",
   163 => x"0402ec05",
   164 => x"0d800b80",
   165 => x"dde40cf6",
   166 => x"8c08f690",
   167 => x"0871882c",
   168 => x"565381ff",
   169 => x"06537373",
   170 => x"25893872",
   171 => x"54820b80",
   172 => x"dde40c71",
   173 => x"882c7281",
   174 => x"ff065355",
   175 => x"7472258d",
   176 => x"387180dd",
   177 => x"e4088407",
   178 => x"80dde40c",
   179 => x"5573842b",
   180 => x"75832b56",
   181 => x"5483f474",
   182 => x"258f3883",
   183 => x"0b0b0b80",
   184 => x"d3d00c82",
   185 => x"985385f3",
   186 => x"04810b0b",
   187 => x"0b80d3d0",
   188 => x"0ca8530b",
   189 => x"0b80d3d0",
   190 => x"0881712b",
   191 => x"ff05f688",
   192 => x"0c747431",
   193 => x"ffb005ff",
   194 => x"1271712c",
   195 => x"ff941970",
   196 => x"9f2a1170",
   197 => x"812c80dd",
   198 => x"e4085255",
   199 => x"51525652",
   200 => x"53517680",
   201 => x"2e853870",
   202 => x"81075170",
   203 => x"f6940c72",
   204 => x"098105f6",
   205 => x"800c7109",
   206 => x"8105f684",
   207 => x"0c029405",
   208 => x"0d040402",
   209 => x"fc050d80",
   210 => x"d9f0519b",
   211 => x"932d0284",
   212 => x"050d0402",
   213 => x"fc050d80",
   214 => x"d3d4519b",
   215 => x"932d0284",
   216 => x"050d0402",
   217 => x"fc050d80",
   218 => x"d8c8519b",
   219 => x"932d0284",
   220 => x"050d0402",
   221 => x"fc050d81",
   222 => x"808051c0",
   223 => x"115170fb",
   224 => x"38028405",
   225 => x"0d047181",
   226 => x"2e098106",
   227 => x"893881c3",
   228 => x"0bec0c87",
   229 => x"9a04830b",
   230 => x"ec0c86f3",
   231 => x"2d820bec",
   232 => x"0c0498d6",
   233 => x"2d80ddcc",
   234 => x"0880d8b8",
   235 => x"0c98d62d",
   236 => x"80ddcc08",
   237 => x"80d7e40c",
   238 => x"98d62d80",
   239 => x"ddcc0880",
   240 => x"db880c98",
   241 => x"d62d80dd",
   242 => x"cc0880d9",
   243 => x"e00c98d6",
   244 => x"2d80ddcc",
   245 => x"0880d4f8",
   246 => x"0c0402fc",
   247 => x"050d84bf",
   248 => x"5186f32d",
   249 => x"ff115170",
   250 => x"8025f638",
   251 => x"0284050d",
   252 => x"0402f405",
   253 => x"0d745372",
   254 => x"70810554",
   255 => x"80f52d52",
   256 => x"71802e89",
   257 => x"38715183",
   258 => x"842d87f7",
   259 => x"04810b80",
   260 => x"ddcc0c02",
   261 => x"8c050d04",
   262 => x"02e8050d",
   263 => x"800b80dd",
   264 => x"f40c800b",
   265 => x"80dbe00c",
   266 => x"80d5c80b",
   267 => x"80f52d51",
   268 => x"70b12e09",
   269 => x"81068d38",
   270 => x"810b80db",
   271 => x"e00c810b",
   272 => x"80ddf40c",
   273 => x"80d5c90b",
   274 => x"80f52d51",
   275 => x"70b12e09",
   276 => x"81069538",
   277 => x"80dbe008",
   278 => x"820780db",
   279 => x"e00c80dd",
   280 => x"f4088207",
   281 => x"80ddf40c",
   282 => x"80d5ca0b",
   283 => x"80f52d51",
   284 => x"70b12e09",
   285 => x"81069538",
   286 => x"80dbe008",
   287 => x"840780db",
   288 => x"e00c80dd",
   289 => x"f4088407",
   290 => x"80ddf40c",
   291 => x"80d5cb0b",
   292 => x"80f52d51",
   293 => x"70b12e09",
   294 => x"81069538",
   295 => x"80dbe008",
   296 => x"880780db",
   297 => x"e00c80dd",
   298 => x"f4088807",
   299 => x"80ddf40c",
   300 => x"80d5cc0b",
   301 => x"80f52d51",
   302 => x"70b12e09",
   303 => x"81069538",
   304 => x"80dbe008",
   305 => x"900780db",
   306 => x"e00c80dd",
   307 => x"f4089007",
   308 => x"80ddf40c",
   309 => x"80d5cd0b",
   310 => x"80f52d51",
   311 => x"70b12e09",
   312 => x"81069538",
   313 => x"80dbe008",
   314 => x"a00780db",
   315 => x"e00c80dd",
   316 => x"f408a007",
   317 => x"80ddf40c",
   318 => x"80d5ce0b",
   319 => x"80f52d51",
   320 => x"70b12e09",
   321 => x"81069d38",
   322 => x"80dbe008",
   323 => x"80c00780",
   324 => x"dbe00c80",
   325 => x"ddf40880",
   326 => x"c00780dd",
   327 => x"f40c810b",
   328 => x"80d5d80c",
   329 => x"80d5cf0b",
   330 => x"80f52dd0",
   331 => x"05517080",
   332 => x"d3f40b81",
   333 => x"b72d80d5",
   334 => x"d00b80f5",
   335 => x"2dd00554",
   336 => x"7380d480",
   337 => x"0b81b72d",
   338 => x"80d5d10b",
   339 => x"80f52dd0",
   340 => x"05557480",
   341 => x"d4980b81",
   342 => x"b72d80d5",
   343 => x"d20b80f5",
   344 => x"2dd00552",
   345 => x"7180d4b0",
   346 => x"0b81b72d",
   347 => x"80d5d30b",
   348 => x"80f52dd0",
   349 => x"05537280",
   350 => x"d4e00b81",
   351 => x"b72d708a",
   352 => x"2b8ff880",
   353 => x"06748b2b",
   354 => x"9ff08006",
   355 => x"7180ddf4",
   356 => x"08070776",
   357 => x"8d2b80ff",
   358 => x"c0800674",
   359 => x"8e2b81ff",
   360 => x"80800671",
   361 => x"73070776",
   362 => x"912b8ff8",
   363 => x"80800671",
   364 => x"077080dd",
   365 => x"f40cfc0c",
   366 => x"52575151",
   367 => x"0298050d",
   368 => x"0402f805",
   369 => x"0d810bec",
   370 => x"0c840bec",
   371 => x"0c80c6b8",
   372 => x"5280dde8",
   373 => x"51bb952d",
   374 => x"80ddcc08",
   375 => x"802e81bd",
   376 => x"3880dec4",
   377 => x"5280dde8",
   378 => x"51be882d",
   379 => x"80ddcc08",
   380 => x"802e81a9",
   381 => x"3880dec4",
   382 => x"0b80f52d",
   383 => x"80d5c80b",
   384 => x"81b72d80",
   385 => x"dec50b80",
   386 => x"f52d80d5",
   387 => x"c90b81b7",
   388 => x"2d80dec6",
   389 => x"0b80f52d",
   390 => x"80d5ca0b",
   391 => x"81b72d80",
   392 => x"dec70b80",
   393 => x"f52d80d5",
   394 => x"cb0b81b7",
   395 => x"2d80dec8",
   396 => x"0b80f52d",
   397 => x"80d5cc0b",
   398 => x"81b72d80",
   399 => x"dec90b80",
   400 => x"f52d80d5",
   401 => x"cd0b81b7",
   402 => x"2d80deca",
   403 => x"0b80f52d",
   404 => x"80d5ce0b",
   405 => x"81b72d80",
   406 => x"decb0b80",
   407 => x"f52d80d5",
   408 => x"cf0b81b7",
   409 => x"2d80decc",
   410 => x"0b80f52d",
   411 => x"80d5d00b",
   412 => x"81b72d80",
   413 => x"decd0b80",
   414 => x"f52d80d5",
   415 => x"d10b81b7",
   416 => x"2d80dece",
   417 => x"0b80f52d",
   418 => x"80d5d20b",
   419 => x"81b72d80",
   420 => x"decf0b80",
   421 => x"f52d80d5",
   422 => x"d30b81b7",
   423 => x"2d88982d",
   424 => x"0288050d",
   425 => x"0402dc05",
   426 => x"0d800b80",
   427 => x"d5dc0854",
   428 => x"5972832e",
   429 => x"a8387283",
   430 => x"24893872",
   431 => x"822e8c38",
   432 => x"8e810472",
   433 => x"842ea838",
   434 => x"8e810480",
   435 => x"ddf408bf",
   436 => x"faff0682",
   437 => x"800780dd",
   438 => x"f40c8e90",
   439 => x"0480ddf4",
   440 => x"08bfffff",
   441 => x"06878007",
   442 => x"80ddf40c",
   443 => x"8e900480",
   444 => x"ddf408bf",
   445 => x"fbff0683",
   446 => x"800780dd",
   447 => x"f40c8e90",
   448 => x"0480ddf4",
   449 => x"08bff9ff",
   450 => x"06818007",
   451 => x"80ddf40c",
   452 => x"80ddf408",
   453 => x"fc0c8184",
   454 => x"0bec0c7a",
   455 => x"5280dde8",
   456 => x"51bb952d",
   457 => x"80ddcc08",
   458 => x"802e819d",
   459 => x"3880ddec",
   460 => x"08548056",
   461 => x"73852e09",
   462 => x"81068a38",
   463 => x"840bec0c",
   464 => x"81538fd1",
   465 => x"0473f80c",
   466 => x"81a40bec",
   467 => x"0c87da2d",
   468 => x"75ff1557",
   469 => x"5875802e",
   470 => x"8b388118",
   471 => x"76812a57",
   472 => x"588ed504",
   473 => x"f7185881",
   474 => x"59807425",
   475 => x"80d738a4",
   476 => x"0bec0c77",
   477 => x"52755184",
   478 => x"a82d80de",
   479 => x"c45280dd",
   480 => x"e851be88",
   481 => x"2d80ddcc",
   482 => x"08802ea0",
   483 => x"3880dec4",
   484 => x"5783fc55",
   485 => x"76708405",
   486 => x"5808e80c",
   487 => x"fc155574",
   488 => x"8025f138",
   489 => x"81a40bec",
   490 => x"0c8fb404",
   491 => x"80ddcc08",
   492 => x"59848054",
   493 => x"80dde851",
   494 => x"bdd82dfc",
   495 => x"80148117",
   496 => x"57548ee9",
   497 => x"04840bec",
   498 => x"0c80ddec",
   499 => x"08f80c78",
   500 => x"537280dd",
   501 => x"cc0c02a4",
   502 => x"050d0402",
   503 => x"f8050d73",
   504 => x"518da52d",
   505 => x"80ddcc08",
   506 => x"5280ddcc",
   507 => x"08802e88",
   508 => x"3880d7f4",
   509 => x"518ffc04",
   510 => x"80d7d051",
   511 => x"9b932d71",
   512 => x"80ddcc0c",
   513 => x"0288050d",
   514 => x"0402f005",
   515 => x"0d800b80",
   516 => x"ddf40c81",
   517 => x"5187862d",
   518 => x"80518786",
   519 => x"2d840bec",
   520 => x"0c98a62d",
   521 => x"94d12d81",
   522 => x"f92d8352",
   523 => x"98892d81",
   524 => x"51858d2d",
   525 => x"ff125271",
   526 => x"8025f138",
   527 => x"80c40bec",
   528 => x"0c80d1a0",
   529 => x"5187f12d",
   530 => x"b1b62d80",
   531 => x"ddcc0880",
   532 => x"2e83e738",
   533 => x"81840bec",
   534 => x"0c80d1b8",
   535 => x"5187f12d",
   536 => x"80ddf408",
   537 => x"bfffff06",
   538 => x"87800770",
   539 => x"80ddf40c",
   540 => x"fc0c80d1",
   541 => x"d0518da5",
   542 => x"2d80ddcc",
   543 => x"08802e80",
   544 => x"df3880d1",
   545 => x"dc518da5",
   546 => x"2d80ddcc",
   547 => x"08802ebd",
   548 => x"3880d1e8",
   549 => x"518da52d",
   550 => x"80ddcc08",
   551 => x"5280ddcc",
   552 => x"08973880",
   553 => x"d1f45187",
   554 => x"f12d80d2",
   555 => x"8c518da5",
   556 => x"2d715187",
   557 => x"862d91d4",
   558 => x"0480d28c",
   559 => x"518da52d",
   560 => x"80518786",
   561 => x"2d805185",
   562 => x"8d2d91d4",
   563 => x"0480d1f4",
   564 => x"5187f12d",
   565 => x"8bc12dfc",
   566 => x"0880ddf4",
   567 => x"0c91e704",
   568 => x"80d1f451",
   569 => x"87f12d84",
   570 => x"0bec0c8f",
   571 => x"db5180c6",
   572 => x"9f2d80dd",
   573 => x"f408fc0c",
   574 => x"80dea408",
   575 => x"882a7081",
   576 => x"06515271",
   577 => x"802e8c38",
   578 => x"80d6d80b",
   579 => x"80ddf80c",
   580 => x"929b0480",
   581 => x"d5e00b80",
   582 => x"ddf80c80",
   583 => x"ddf80851",
   584 => x"9b932d80",
   585 => x"5187a22d",
   586 => x"830b80de",
   587 => x"b80c98df",
   588 => x"2d805185",
   589 => x"8d2d98f3",
   590 => x"2d94dd2d",
   591 => x"9ba62d80",
   592 => x"d3f40b80",
   593 => x"f52d80d4",
   594 => x"800b80f5",
   595 => x"2d718a2b",
   596 => x"718b2b07",
   597 => x"80d4980b",
   598 => x"80f52d70",
   599 => x"8d2b7207",
   600 => x"80d4b00b",
   601 => x"80f52d70",
   602 => x"8e2b7207",
   603 => x"80d4e00b",
   604 => x"80f52d70",
   605 => x"912b7207",
   606 => x"7080ddf4",
   607 => x"0c80dbe0",
   608 => x"08708106",
   609 => x"54525354",
   610 => x"52545253",
   611 => x"54555371",
   612 => x"802e8838",
   613 => x"73810780",
   614 => x"ddf40c72",
   615 => x"812a7081",
   616 => x"06515271",
   617 => x"802e8b38",
   618 => x"80ddf408",
   619 => x"820780dd",
   620 => x"f40c7282",
   621 => x"2a708106",
   622 => x"51527180",
   623 => x"2e8b3880",
   624 => x"ddf40884",
   625 => x"0780ddf4",
   626 => x"0c72832a",
   627 => x"70810651",
   628 => x"5271802e",
   629 => x"8b3880dd",
   630 => x"f4088807",
   631 => x"80ddf40c",
   632 => x"72842a70",
   633 => x"81065152",
   634 => x"71802e8b",
   635 => x"3880ddf4",
   636 => x"08900780",
   637 => x"ddf40c72",
   638 => x"852a7081",
   639 => x"06515271",
   640 => x"802e8b38",
   641 => x"80ddf408",
   642 => x"a00780dd",
   643 => x"f40c80d5",
   644 => x"d808812e",
   645 => x"0981068c",
   646 => x"3880ddf4",
   647 => x"0880c007",
   648 => x"80ddf40c",
   649 => x"80ddf408",
   650 => x"fc0c8652",
   651 => x"80ddcc08",
   652 => x"83388452",
   653 => x"71ec0c92",
   654 => x"b904800b",
   655 => x"80ddcc0c",
   656 => x"0290050d",
   657 => x"0471980c",
   658 => x"04ffb008",
   659 => x"80ddcc0c",
   660 => x"04810bff",
   661 => x"b00c0480",
   662 => x"0bffb00c",
   663 => x"0402f405",
   664 => x"0d95eb04",
   665 => x"80ddcc08",
   666 => x"81f02e09",
   667 => x"81068a38",
   668 => x"810b80db",
   669 => x"d80c95eb",
   670 => x"0480ddcc",
   671 => x"0881e02e",
   672 => x"0981068a",
   673 => x"38810b80",
   674 => x"dbdc0c95",
   675 => x"eb0480dd",
   676 => x"cc085280",
   677 => x"dbdc0880",
   678 => x"2e893880",
   679 => x"ddcc0881",
   680 => x"80055271",
   681 => x"842c728f",
   682 => x"06535380",
   683 => x"dbd80880",
   684 => x"2e9a3872",
   685 => x"842980db",
   686 => x"98057213",
   687 => x"81712b70",
   688 => x"09730806",
   689 => x"730c5153",
   690 => x"5395df04",
   691 => x"72842980",
   692 => x"db980572",
   693 => x"1383712b",
   694 => x"72080772",
   695 => x"0c535380",
   696 => x"0b80dbdc",
   697 => x"0c800b80",
   698 => x"dbd80c80",
   699 => x"ddfc5196",
   700 => x"f22d80dd",
   701 => x"cc08ff24",
   702 => x"feea3880",
   703 => x"0b80ddcc",
   704 => x"0c028c05",
   705 => x"0d0402f8",
   706 => x"050d80db",
   707 => x"98528f51",
   708 => x"80727084",
   709 => x"05540cff",
   710 => x"11517080",
   711 => x"25f23802",
   712 => x"88050d04",
   713 => x"02f0050d",
   714 => x"755194d7",
   715 => x"2d70822c",
   716 => x"fc0680db",
   717 => x"98117210",
   718 => x"9e067108",
   719 => x"70722a70",
   720 => x"83068274",
   721 => x"2b700974",
   722 => x"06760c54",
   723 => x"51565753",
   724 => x"515394d1",
   725 => x"2d7180dd",
   726 => x"cc0c0290",
   727 => x"050d0402",
   728 => x"fc050d72",
   729 => x"5180710c",
   730 => x"800b8412",
   731 => x"0c028405",
   732 => x"0d0402f0",
   733 => x"050d7570",
   734 => x"08841208",
   735 => x"535353ff",
   736 => x"5471712e",
   737 => x"a83894d7",
   738 => x"2d841308",
   739 => x"70842914",
   740 => x"88117008",
   741 => x"7081ff06",
   742 => x"84180881",
   743 => x"11870684",
   744 => x"1a0c5351",
   745 => x"55515151",
   746 => x"94d12d71",
   747 => x"547380dd",
   748 => x"cc0c0290",
   749 => x"050d0402",
   750 => x"f4050d94",
   751 => x"d72de008",
   752 => x"708b2a70",
   753 => x"81065152",
   754 => x"5370802e",
   755 => x"a13880dd",
   756 => x"fc087084",
   757 => x"2980de84",
   758 => x"057481ff",
   759 => x"06710c51",
   760 => x"5180ddfc",
   761 => x"08811187",
   762 => x"0680ddfc",
   763 => x"0c51728c",
   764 => x"2c83ff06",
   765 => x"80dea40c",
   766 => x"800b80de",
   767 => x"a80c94c9",
   768 => x"2d94d12d",
   769 => x"028c050d",
   770 => x"0402fc05",
   771 => x"0d94d72d",
   772 => x"810b80de",
   773 => x"a80c94d1",
   774 => x"2d80dea8",
   775 => x"085170f9",
   776 => x"38028405",
   777 => x"0d0402fc",
   778 => x"050d80dd",
   779 => x"fc5196df",
   780 => x"2d96862d",
   781 => x"97b75194",
   782 => x"c52d0284",
   783 => x"050d0402",
   784 => x"fc050d8f",
   785 => x"cf5186f3",
   786 => x"2dff1151",
   787 => x"708025f6",
   788 => x"38028405",
   789 => x"0d0480de",
   790 => x"b00880dd",
   791 => x"cc0c0402",
   792 => x"fc050d81",
   793 => x"0b80dc8c",
   794 => x"0c815185",
   795 => x"8d2d0284",
   796 => x"050d0402",
   797 => x"f8050d98",
   798 => x"fd0494dd",
   799 => x"2d80da51",
   800 => x"96a42d80",
   801 => x"ddcc0881",
   802 => x"065271ee",
   803 => x"3880dc88",
   804 => x"085196a4",
   805 => x"2d80ddcc",
   806 => x"08810652",
   807 => x"71dc3883",
   808 => x"5196a42d",
   809 => x"80ddcc08",
   810 => x"81065271",
   811 => x"cd387180",
   812 => x"dc8c0c71",
   813 => x"51858d2d",
   814 => x"0288050d",
   815 => x"0402ec05",
   816 => x"0d765480",
   817 => x"52870b88",
   818 => x"1580f52d",
   819 => x"56537472",
   820 => x"248338a0",
   821 => x"53725183",
   822 => x"842d8112",
   823 => x"8b1580f5",
   824 => x"2d545272",
   825 => x"7225de38",
   826 => x"0294050d",
   827 => x"0402f005",
   828 => x"0d80deb0",
   829 => x"085481f9",
   830 => x"2d800b80",
   831 => x"deb40c73",
   832 => x"08802e81",
   833 => x"8938820b",
   834 => x"80dde00c",
   835 => x"80deb408",
   836 => x"8f0680dd",
   837 => x"dc0c7308",
   838 => x"5271832e",
   839 => x"96387183",
   840 => x"26893871",
   841 => x"812eb038",
   842 => x"9af70471",
   843 => x"852ea038",
   844 => x"9af70488",
   845 => x"1480f52d",
   846 => x"84150880",
   847 => x"d2985354",
   848 => x"5287f12d",
   849 => x"71842913",
   850 => x"70085252",
   851 => x"9afb0473",
   852 => x"5199bd2d",
   853 => x"9af70480",
   854 => x"dbe00888",
   855 => x"15082c70",
   856 => x"81065152",
   857 => x"71802e88",
   858 => x"3880d29c",
   859 => x"519af404",
   860 => x"80d2a051",
   861 => x"87f12d84",
   862 => x"14085187",
   863 => x"f12d80de",
   864 => x"b4088105",
   865 => x"80deb40c",
   866 => x"8c145499",
   867 => x"ff040290",
   868 => x"050d0471",
   869 => x"80deb00c",
   870 => x"99ed2d80",
   871 => x"deb408ff",
   872 => x"0580deb8",
   873 => x"0c0402e8",
   874 => x"050d80de",
   875 => x"b00880de",
   876 => x"bc085755",
   877 => x"835196a4",
   878 => x"2d80ddcc",
   879 => x"08830652",
   880 => x"71802ea5",
   881 => x"389bcb04",
   882 => x"94dd2d83",
   883 => x"5196a42d",
   884 => x"80ddcc08",
   885 => x"81065271",
   886 => x"ef3880dc",
   887 => x"8c088132",
   888 => x"7080dc8c",
   889 => x"0c51858d",
   890 => x"2d800b80",
   891 => x"deac0c8c",
   892 => x"5196a42d",
   893 => x"80ddcc08",
   894 => x"812a7081",
   895 => x"06515271",
   896 => x"802e80d1",
   897 => x"3880dbe4",
   898 => x"0880dbf8",
   899 => x"0880dbe4",
   900 => x"0c80dbf8",
   901 => x"0c80dbe8",
   902 => x"0880dbfc",
   903 => x"0880dbe8",
   904 => x"0c80dbfc",
   905 => x"0c80dbec",
   906 => x"0880dc80",
   907 => x"0880dbec",
   908 => x"0c80dc80",
   909 => x"0c80dbf0",
   910 => x"0880dc84",
   911 => x"0880dbf0",
   912 => x"0c80dc84",
   913 => x"0c80dbf4",
   914 => x"0880dc88",
   915 => x"0880dbf4",
   916 => x"0c80dc88",
   917 => x"0c80dea4",
   918 => x"08a00652",
   919 => x"80722596",
   920 => x"3898bf2d",
   921 => x"94dd2d80",
   922 => x"dc8c0881",
   923 => x"327080dc",
   924 => x"8c0c5185",
   925 => x"8d2d80dc",
   926 => x"8c0883a4",
   927 => x"3880dbf8",
   928 => x"085196a4",
   929 => x"2d80ddcc",
   930 => x"08802e8b",
   931 => x"3880deac",
   932 => x"08810780",
   933 => x"deac0c80",
   934 => x"dbfc0851",
   935 => x"96a42d80",
   936 => x"ddcc0880",
   937 => x"2e8b3880",
   938 => x"deac0882",
   939 => x"0780deac",
   940 => x"0c80dc80",
   941 => x"085196a4",
   942 => x"2d80ddcc",
   943 => x"08802e8b",
   944 => x"3880deac",
   945 => x"08840780",
   946 => x"deac0c80",
   947 => x"dc840851",
   948 => x"96a42d80",
   949 => x"ddcc0880",
   950 => x"2e8b3880",
   951 => x"deac0888",
   952 => x"0780deac",
   953 => x"0c80dc88",
   954 => x"085196a4",
   955 => x"2d80ddcc",
   956 => x"08802e8b",
   957 => x"3880deac",
   958 => x"08900780",
   959 => x"deac0c80",
   960 => x"dbe40851",
   961 => x"96a42d80",
   962 => x"ddcc0880",
   963 => x"2e8c3880",
   964 => x"deac0882",
   965 => x"800780de",
   966 => x"ac0c80db",
   967 => x"e8085196",
   968 => x"a42d80dd",
   969 => x"cc08802e",
   970 => x"8c3880de",
   971 => x"ac088480",
   972 => x"0780deac",
   973 => x"0c80dbec",
   974 => x"085196a4",
   975 => x"2d80ddcc",
   976 => x"08802e8c",
   977 => x"3880deac",
   978 => x"08888007",
   979 => x"80deac0c",
   980 => x"80dbf008",
   981 => x"5196a42d",
   982 => x"80ddcc08",
   983 => x"802e8c38",
   984 => x"80deac08",
   985 => x"90800780",
   986 => x"deac0c80",
   987 => x"dbf40851",
   988 => x"96a42d80",
   989 => x"ddcc0880",
   990 => x"2e8c3880",
   991 => x"deac08a0",
   992 => x"800780de",
   993 => x"ac0c9451",
   994 => x"96a42d80",
   995 => x"ddcc0852",
   996 => x"915196a4",
   997 => x"2d7180dd",
   998 => x"cc080652",
   999 => x"80e65196",
  1000 => x"a42d7180",
  1001 => x"ddcc0806",
  1002 => x"5271802e",
  1003 => x"8d3880de",
  1004 => x"ac088480",
  1005 => x"800780de",
  1006 => x"ac0c80fe",
  1007 => x"5196a42d",
  1008 => x"80ddcc08",
  1009 => x"52875196",
  1010 => x"a42d7180",
  1011 => x"ddcc0807",
  1012 => x"5271802e",
  1013 => x"8d3880de",
  1014 => x"ac088880",
  1015 => x"800780de",
  1016 => x"ac0c80de",
  1017 => x"ac08ed0c",
  1018 => x"8a5196a4",
  1019 => x"2d80ddcc",
  1020 => x"08812a70",
  1021 => x"81065152",
  1022 => x"71802e89",
  1023 => x"8e38a084",
  1024 => x"0494dd2d",
  1025 => x"8a5196a4",
  1026 => x"2d80ddcc",
  1027 => x"08810652",
  1028 => x"71ef3880",
  1029 => x"d5d80881",
  1030 => x"3280d5d8",
  1031 => x"0ca98b04",
  1032 => x"945196a4",
  1033 => x"2d80ddcc",
  1034 => x"08529151",
  1035 => x"96a42d71",
  1036 => x"80ddcc08",
  1037 => x"065280e6",
  1038 => x"5196a42d",
  1039 => x"7180ddcc",
  1040 => x"08065271",
  1041 => x"802e8d38",
  1042 => x"80deac08",
  1043 => x"84808007",
  1044 => x"80deac0c",
  1045 => x"80fe5196",
  1046 => x"a42d80dd",
  1047 => x"cc085287",
  1048 => x"5196a42d",
  1049 => x"7180ddcc",
  1050 => x"08075271",
  1051 => x"802e8d38",
  1052 => x"80deac08",
  1053 => x"88808007",
  1054 => x"80deac0c",
  1055 => x"8a5196a4",
  1056 => x"2d80ddcc",
  1057 => x"08812a70",
  1058 => x"81065152",
  1059 => x"71802ea0",
  1060 => x"38a19704",
  1061 => x"94dd2d8a",
  1062 => x"5196a42d",
  1063 => x"80ddcc08",
  1064 => x"81065271",
  1065 => x"ef3880d5",
  1066 => x"d8088132",
  1067 => x"80d5d80c",
  1068 => x"80deac08",
  1069 => x"ed0c81f5",
  1070 => x"5196a42d",
  1071 => x"80ddcc08",
  1072 => x"812a7081",
  1073 => x"06515271",
  1074 => x"a43880db",
  1075 => x"f8085196",
  1076 => x"a42d80dd",
  1077 => x"cc08812a",
  1078 => x"70810651",
  1079 => x"52718e38",
  1080 => x"80dea408",
  1081 => x"81065280",
  1082 => x"722580c2",
  1083 => x"3880dea4",
  1084 => x"08810652",
  1085 => x"80722584",
  1086 => x"3898bf2d",
  1087 => x"80deb808",
  1088 => x"5271802e",
  1089 => x"8a38ff12",
  1090 => x"80deb80c",
  1091 => x"a2ae0480",
  1092 => x"deb40810",
  1093 => x"80deb408",
  1094 => x"05708429",
  1095 => x"16515288",
  1096 => x"1208802e",
  1097 => x"8938ff51",
  1098 => x"88120852",
  1099 => x"712d81f2",
  1100 => x"5196a42d",
  1101 => x"80ddcc08",
  1102 => x"812a7081",
  1103 => x"06515271",
  1104 => x"a43880db",
  1105 => x"fc085196",
  1106 => x"a42d80dd",
  1107 => x"cc08812a",
  1108 => x"70810651",
  1109 => x"52718e38",
  1110 => x"80dea408",
  1111 => x"82065280",
  1112 => x"722580c3",
  1113 => x"3880dea4",
  1114 => x"08820652",
  1115 => x"80722584",
  1116 => x"3898bf2d",
  1117 => x"80deb408",
  1118 => x"ff1180de",
  1119 => x"b8085653",
  1120 => x"53737225",
  1121 => x"8a388114",
  1122 => x"80deb80c",
  1123 => x"a3a70472",
  1124 => x"10137084",
  1125 => x"29165152",
  1126 => x"88120880",
  1127 => x"2e8938fe",
  1128 => x"51881208",
  1129 => x"52712d81",
  1130 => x"fd5196a4",
  1131 => x"2d80ddcc",
  1132 => x"08812a70",
  1133 => x"81065152",
  1134 => x"71ba3880",
  1135 => x"dc800851",
  1136 => x"96a42d80",
  1137 => x"ddcc0881",
  1138 => x"2a708106",
  1139 => x"515271a4",
  1140 => x"3880dea4",
  1141 => x"08840652",
  1142 => x"71802498",
  1143 => x"3881eb51",
  1144 => x"96a42d80",
  1145 => x"ddcc0881",
  1146 => x"2a708106",
  1147 => x"51527180",
  1148 => x"2e80c038",
  1149 => x"80dea408",
  1150 => x"84065280",
  1151 => x"72258438",
  1152 => x"98bf2d80",
  1153 => x"deb80880",
  1154 => x"2e8a3880",
  1155 => x"0b80deb8",
  1156 => x"0ca4b304",
  1157 => x"80deb408",
  1158 => x"1080deb4",
  1159 => x"08057084",
  1160 => x"29165152",
  1161 => x"88120880",
  1162 => x"2e8938fd",
  1163 => x"51881208",
  1164 => x"52712d81",
  1165 => x"fa5196a4",
  1166 => x"2d80ddcc",
  1167 => x"08812a70",
  1168 => x"81065152",
  1169 => x"71ba3880",
  1170 => x"dc840851",
  1171 => x"96a42d80",
  1172 => x"ddcc0881",
  1173 => x"2a708106",
  1174 => x"515271a4",
  1175 => x"3880dea4",
  1176 => x"08880652",
  1177 => x"71802498",
  1178 => x"3881f451",
  1179 => x"96a42d80",
  1180 => x"ddcc0881",
  1181 => x"2a708106",
  1182 => x"51527180",
  1183 => x"2e80c038",
  1184 => x"80dea408",
  1185 => x"88065280",
  1186 => x"72258438",
  1187 => x"98bf2d80",
  1188 => x"deb408ff",
  1189 => x"11545280",
  1190 => x"deb80873",
  1191 => x"25893872",
  1192 => x"80deb80c",
  1193 => x"a5bf0471",
  1194 => x"10127084",
  1195 => x"29165152",
  1196 => x"88120880",
  1197 => x"2e8938fc",
  1198 => x"51881208",
  1199 => x"52712d80",
  1200 => x"deb80870",
  1201 => x"53547380",
  1202 => x"2e8a388c",
  1203 => x"15ff1555",
  1204 => x"55a5c604",
  1205 => x"820b80dd",
  1206 => x"e00c718f",
  1207 => x"0680dddc",
  1208 => x"0c81eb51",
  1209 => x"96a42d80",
  1210 => x"ddcc0881",
  1211 => x"2a708106",
  1212 => x"51527180",
  1213 => x"2ead3874",
  1214 => x"08852e09",
  1215 => x"8106a438",
  1216 => x"881580f5",
  1217 => x"2dff0552",
  1218 => x"71881681",
  1219 => x"b72d7198",
  1220 => x"2b527180",
  1221 => x"25883880",
  1222 => x"0b881681",
  1223 => x"b72d7451",
  1224 => x"99bd2d81",
  1225 => x"f45196a4",
  1226 => x"2d80ddcc",
  1227 => x"08812a70",
  1228 => x"81065152",
  1229 => x"71802eb3",
  1230 => x"38740885",
  1231 => x"2e098106",
  1232 => x"aa388815",
  1233 => x"80f52d81",
  1234 => x"05527188",
  1235 => x"1681b72d",
  1236 => x"7181ff06",
  1237 => x"8b1680f5",
  1238 => x"2d545272",
  1239 => x"72278738",
  1240 => x"72881681",
  1241 => x"b72d7451",
  1242 => x"99bd2d80",
  1243 => x"da5196a4",
  1244 => x"2d80ddcc",
  1245 => x"08812a70",
  1246 => x"81065152",
  1247 => x"718e3880",
  1248 => x"dea40890",
  1249 => x"06528072",
  1250 => x"2581bc38",
  1251 => x"80deb008",
  1252 => x"80dea408",
  1253 => x"90065353",
  1254 => x"80722584",
  1255 => x"3898bf2d",
  1256 => x"80deb808",
  1257 => x"5473802e",
  1258 => x"8a388c13",
  1259 => x"ff155553",
  1260 => x"a7a50472",
  1261 => x"08527182",
  1262 => x"2ea63871",
  1263 => x"82268938",
  1264 => x"71812eaa",
  1265 => x"38a8c704",
  1266 => x"71832eb4",
  1267 => x"3871842e",
  1268 => x"09810680",
  1269 => x"f2388813",
  1270 => x"08519b93",
  1271 => x"2da8c704",
  1272 => x"80deb808",
  1273 => x"51881308",
  1274 => x"52712da8",
  1275 => x"c704810b",
  1276 => x"8814082b",
  1277 => x"80dbe008",
  1278 => x"3280dbe0",
  1279 => x"0ca89b04",
  1280 => x"881380f5",
  1281 => x"2d81058b",
  1282 => x"1480f52d",
  1283 => x"53547174",
  1284 => x"24833880",
  1285 => x"54738814",
  1286 => x"81b72d99",
  1287 => x"ed2da8c7",
  1288 => x"04750880",
  1289 => x"2ea43875",
  1290 => x"085196a4",
  1291 => x"2d80ddcc",
  1292 => x"08810652",
  1293 => x"71802e8c",
  1294 => x"3880deb8",
  1295 => x"08518416",
  1296 => x"0852712d",
  1297 => x"88165675",
  1298 => x"d8388054",
  1299 => x"800b80dd",
  1300 => x"e00c738f",
  1301 => x"0680dddc",
  1302 => x"0ca05273",
  1303 => x"80deb808",
  1304 => x"2e098106",
  1305 => x"993880de",
  1306 => x"b408ff05",
  1307 => x"74327009",
  1308 => x"81057072",
  1309 => x"079f2a91",
  1310 => x"71315151",
  1311 => x"53537151",
  1312 => x"83842d81",
  1313 => x"14548e74",
  1314 => x"25c23880",
  1315 => x"dc8c0880",
  1316 => x"ddcc0c02",
  1317 => x"98050d04",
  1318 => x"02f4050d",
  1319 => x"d45281ff",
  1320 => x"720c7108",
  1321 => x"5381ff72",
  1322 => x"0c72882b",
  1323 => x"83fe8006",
  1324 => x"72087081",
  1325 => x"ff065152",
  1326 => x"5381ff72",
  1327 => x"0c727107",
  1328 => x"882b7208",
  1329 => x"7081ff06",
  1330 => x"51525381",
  1331 => x"ff720c72",
  1332 => x"7107882b",
  1333 => x"72087081",
  1334 => x"ff067207",
  1335 => x"80ddcc0c",
  1336 => x"5253028c",
  1337 => x"050d0402",
  1338 => x"f4050d74",
  1339 => x"767181ff",
  1340 => x"06d40c53",
  1341 => x"5380dec0",
  1342 => x"08853871",
  1343 => x"892b5271",
  1344 => x"982ad40c",
  1345 => x"71902a70",
  1346 => x"81ff06d4",
  1347 => x"0c517188",
  1348 => x"2a7081ff",
  1349 => x"06d40c51",
  1350 => x"7181ff06",
  1351 => x"d40c7290",
  1352 => x"2a7081ff",
  1353 => x"06d40c51",
  1354 => x"d4087081",
  1355 => x"ff065151",
  1356 => x"82b8bf52",
  1357 => x"7081ff2e",
  1358 => x"09810694",
  1359 => x"3881ff0b",
  1360 => x"d40cd408",
  1361 => x"7081ff06",
  1362 => x"ff145451",
  1363 => x"5171e538",
  1364 => x"7080ddcc",
  1365 => x"0c028c05",
  1366 => x"0d0402fc",
  1367 => x"050d81c7",
  1368 => x"5181ff0b",
  1369 => x"d40cff11",
  1370 => x"51708025",
  1371 => x"f4380284",
  1372 => x"050d0402",
  1373 => x"f4050d81",
  1374 => x"ff0bd40c",
  1375 => x"93538052",
  1376 => x"87fc80c1",
  1377 => x"51a9e72d",
  1378 => x"80ddcc08",
  1379 => x"8b3881ff",
  1380 => x"0bd40c81",
  1381 => x"53aba104",
  1382 => x"aada2dff",
  1383 => x"135372de",
  1384 => x"387280dd",
  1385 => x"cc0c028c",
  1386 => x"050d0402",
  1387 => x"ec050d81",
  1388 => x"0b80dec0",
  1389 => x"0c8454d0",
  1390 => x"08708f2a",
  1391 => x"70810651",
  1392 => x"515372f3",
  1393 => x"3872d00c",
  1394 => x"aada2d80",
  1395 => x"d2a45187",
  1396 => x"f12dd008",
  1397 => x"708f2a70",
  1398 => x"81065151",
  1399 => x"5372f338",
  1400 => x"810bd00c",
  1401 => x"b1538052",
  1402 => x"84d480c0",
  1403 => x"51a9e72d",
  1404 => x"80ddcc08",
  1405 => x"812e9338",
  1406 => x"72822ebf",
  1407 => x"38ff1353",
  1408 => x"72e438ff",
  1409 => x"145473ff",
  1410 => x"ae38aada",
  1411 => x"2d83aa52",
  1412 => x"849c80c8",
  1413 => x"51a9e72d",
  1414 => x"80ddcc08",
  1415 => x"812e0981",
  1416 => x"069338a9",
  1417 => x"982d80dd",
  1418 => x"cc0883ff",
  1419 => x"ff065372",
  1420 => x"83aa2e9f",
  1421 => x"38aaf32d",
  1422 => x"acce0480",
  1423 => x"d2b05187",
  1424 => x"f12d8053",
  1425 => x"aea30480",
  1426 => x"d2c85187",
  1427 => x"f12d8054",
  1428 => x"adf40481",
  1429 => x"ff0bd40c",
  1430 => x"b154aada",
  1431 => x"2d8fcf53",
  1432 => x"805287fc",
  1433 => x"80f751a9",
  1434 => x"e72d80dd",
  1435 => x"cc085580",
  1436 => x"ddcc0881",
  1437 => x"2e098106",
  1438 => x"9c3881ff",
  1439 => x"0bd40c82",
  1440 => x"0a52849c",
  1441 => x"80e951a9",
  1442 => x"e72d80dd",
  1443 => x"cc08802e",
  1444 => x"8d38aada",
  1445 => x"2dff1353",
  1446 => x"72c638ad",
  1447 => x"e70481ff",
  1448 => x"0bd40c80",
  1449 => x"ddcc0852",
  1450 => x"87fc80fa",
  1451 => x"51a9e72d",
  1452 => x"80ddcc08",
  1453 => x"b23881ff",
  1454 => x"0bd40cd4",
  1455 => x"085381ff",
  1456 => x"0bd40c81",
  1457 => x"ff0bd40c",
  1458 => x"81ff0bd4",
  1459 => x"0c81ff0b",
  1460 => x"d40c7286",
  1461 => x"2a708106",
  1462 => x"76565153",
  1463 => x"72963880",
  1464 => x"ddcc0854",
  1465 => x"adf40473",
  1466 => x"822efedb",
  1467 => x"38ff1454",
  1468 => x"73fee738",
  1469 => x"7380dec0",
  1470 => x"0c738b38",
  1471 => x"815287fc",
  1472 => x"80d051a9",
  1473 => x"e72d81ff",
  1474 => x"0bd40cd0",
  1475 => x"08708f2a",
  1476 => x"70810651",
  1477 => x"515372f3",
  1478 => x"3872d00c",
  1479 => x"81ff0bd4",
  1480 => x"0c815372",
  1481 => x"80ddcc0c",
  1482 => x"0294050d",
  1483 => x"0402e805",
  1484 => x"0d785580",
  1485 => x"5681ff0b",
  1486 => x"d40cd008",
  1487 => x"708f2a70",
  1488 => x"81065151",
  1489 => x"5372f338",
  1490 => x"82810bd0",
  1491 => x"0c81ff0b",
  1492 => x"d40c7752",
  1493 => x"87fc80d1",
  1494 => x"51a9e72d",
  1495 => x"80dbc6df",
  1496 => x"5480ddcc",
  1497 => x"08802e8b",
  1498 => x"3880d2e8",
  1499 => x"5187f12d",
  1500 => x"afc70481",
  1501 => x"ff0bd40c",
  1502 => x"d4087081",
  1503 => x"ff065153",
  1504 => x"7281fe2e",
  1505 => x"0981069e",
  1506 => x"3880ff53",
  1507 => x"a9982d80",
  1508 => x"ddcc0875",
  1509 => x"70840557",
  1510 => x"0cff1353",
  1511 => x"728025ec",
  1512 => x"388156af",
  1513 => x"ac04ff14",
  1514 => x"5473c838",
  1515 => x"81ff0bd4",
  1516 => x"0c81ff0b",
  1517 => x"d40cd008",
  1518 => x"708f2a70",
  1519 => x"81065151",
  1520 => x"5372f338",
  1521 => x"72d00c75",
  1522 => x"80ddcc0c",
  1523 => x"0298050d",
  1524 => x"0402e805",
  1525 => x"0d77797b",
  1526 => x"58555580",
  1527 => x"53727625",
  1528 => x"a3387470",
  1529 => x"81055680",
  1530 => x"f52d7470",
  1531 => x"81055680",
  1532 => x"f52d5252",
  1533 => x"71712e86",
  1534 => x"388151b0",
  1535 => x"86048113",
  1536 => x"53afdd04",
  1537 => x"80517080",
  1538 => x"ddcc0c02",
  1539 => x"98050d04",
  1540 => x"02ec050d",
  1541 => x"76557480",
  1542 => x"2e80c238",
  1543 => x"9a1580e0",
  1544 => x"2d51bee2",
  1545 => x"2d80ddcc",
  1546 => x"0880ddcc",
  1547 => x"0880e6f8",
  1548 => x"0c80ddcc",
  1549 => x"08545480",
  1550 => x"e6d40880",
  1551 => x"2e9a3894",
  1552 => x"1580e02d",
  1553 => x"51bee22d",
  1554 => x"80ddcc08",
  1555 => x"902b83ff",
  1556 => x"f00a0670",
  1557 => x"75075153",
  1558 => x"7280e6f8",
  1559 => x"0c80e6f8",
  1560 => x"08537280",
  1561 => x"2e9d3880",
  1562 => x"e6cc08fe",
  1563 => x"14712980",
  1564 => x"e6e00805",
  1565 => x"80e6fc0c",
  1566 => x"70842b80",
  1567 => x"e6d80c54",
  1568 => x"b1b10480",
  1569 => x"e6e40880",
  1570 => x"e6f80c80",
  1571 => x"e6e80880",
  1572 => x"e6fc0c80",
  1573 => x"e6d40880",
  1574 => x"2e8b3880",
  1575 => x"e6cc0884",
  1576 => x"2b53b1ac",
  1577 => x"0480e6ec",
  1578 => x"08842b53",
  1579 => x"7280e6d8",
  1580 => x"0c029405",
  1581 => x"0d0402d8",
  1582 => x"050d800b",
  1583 => x"80e6d40c",
  1584 => x"8454abab",
  1585 => x"2d80ddcc",
  1586 => x"08802e97",
  1587 => x"3880dec4",
  1588 => x"528051ae",
  1589 => x"ad2d80dd",
  1590 => x"cc08802e",
  1591 => x"8638fe54",
  1592 => x"b1eb04ff",
  1593 => x"14547380",
  1594 => x"24d83873",
  1595 => x"8d3880d2",
  1596 => x"f85187f1",
  1597 => x"2d7355b7",
  1598 => x"c0048056",
  1599 => x"810b80e7",
  1600 => x"800c8853",
  1601 => x"80d38c52",
  1602 => x"80defa51",
  1603 => x"afd12d80",
  1604 => x"ddcc0876",
  1605 => x"2e098106",
  1606 => x"893880dd",
  1607 => x"cc0880e7",
  1608 => x"800c8853",
  1609 => x"80d39852",
  1610 => x"80df9651",
  1611 => x"afd12d80",
  1612 => x"ddcc0889",
  1613 => x"3880ddcc",
  1614 => x"0880e780",
  1615 => x"0c80e780",
  1616 => x"08802e81",
  1617 => x"813880e2",
  1618 => x"8a0b80f5",
  1619 => x"2d80e28b",
  1620 => x"0b80f52d",
  1621 => x"71982b71",
  1622 => x"902b0780",
  1623 => x"e28c0b80",
  1624 => x"f52d7088",
  1625 => x"2b720780",
  1626 => x"e28d0b80",
  1627 => x"f52d7107",
  1628 => x"80e2c20b",
  1629 => x"80f52d80",
  1630 => x"e2c30b80",
  1631 => x"f52d7188",
  1632 => x"2b07535f",
  1633 => x"54525a56",
  1634 => x"57557381",
  1635 => x"abaa2e09",
  1636 => x"81068e38",
  1637 => x"7551beb1",
  1638 => x"2d80ddcc",
  1639 => x"0856b3af",
  1640 => x"047382d4",
  1641 => x"d52e8838",
  1642 => x"80d3a451",
  1643 => x"b3fb0480",
  1644 => x"dec45275",
  1645 => x"51aead2d",
  1646 => x"80ddcc08",
  1647 => x"5580ddcc",
  1648 => x"08802e83",
  1649 => x"fb388853",
  1650 => x"80d39852",
  1651 => x"80df9651",
  1652 => x"afd12d80",
  1653 => x"ddcc088a",
  1654 => x"38810b80",
  1655 => x"e6d40cb4",
  1656 => x"81048853",
  1657 => x"80d38c52",
  1658 => x"80defa51",
  1659 => x"afd12d80",
  1660 => x"ddcc0880",
  1661 => x"2e8b3880",
  1662 => x"d3b85187",
  1663 => x"f12db4e0",
  1664 => x"0480e2c2",
  1665 => x"0b80f52d",
  1666 => x"547380d5",
  1667 => x"2e098106",
  1668 => x"80ce3880",
  1669 => x"e2c30b80",
  1670 => x"f52d5473",
  1671 => x"81aa2e09",
  1672 => x"8106bd38",
  1673 => x"800b80de",
  1674 => x"c40b80f5",
  1675 => x"2d565474",
  1676 => x"81e92e83",
  1677 => x"38815474",
  1678 => x"81eb2e8c",
  1679 => x"38805573",
  1680 => x"752e0981",
  1681 => x"0682f938",
  1682 => x"80decf0b",
  1683 => x"80f52d55",
  1684 => x"748e3880",
  1685 => x"ded00b80",
  1686 => x"f52d5473",
  1687 => x"822e8638",
  1688 => x"8055b7c0",
  1689 => x"0480ded1",
  1690 => x"0b80f52d",
  1691 => x"7080e6cc",
  1692 => x"0cff0580",
  1693 => x"e6d00c80",
  1694 => x"ded20b80",
  1695 => x"f52d80de",
  1696 => x"d30b80f5",
  1697 => x"2d587605",
  1698 => x"77828029",
  1699 => x"057080e6",
  1700 => x"dc0c80de",
  1701 => x"d40b80f5",
  1702 => x"2d7080e6",
  1703 => x"f00c80e6",
  1704 => x"d4085957",
  1705 => x"5876802e",
  1706 => x"81b73888",
  1707 => x"5380d398",
  1708 => x"5280df96",
  1709 => x"51afd12d",
  1710 => x"80ddcc08",
  1711 => x"82823880",
  1712 => x"e6cc0870",
  1713 => x"842b80e6",
  1714 => x"d80c7080",
  1715 => x"e6ec0c80",
  1716 => x"dee90b80",
  1717 => x"f52d80de",
  1718 => x"e80b80f5",
  1719 => x"2d718280",
  1720 => x"290580de",
  1721 => x"ea0b80f5",
  1722 => x"2d708480",
  1723 => x"80291280",
  1724 => x"deeb0b80",
  1725 => x"f52d7081",
  1726 => x"800a2912",
  1727 => x"7080e6f4",
  1728 => x"0c80e6f0",
  1729 => x"08712980",
  1730 => x"e6dc0805",
  1731 => x"7080e6e0",
  1732 => x"0c80def1",
  1733 => x"0b80f52d",
  1734 => x"80def00b",
  1735 => x"80f52d71",
  1736 => x"82802905",
  1737 => x"80def20b",
  1738 => x"80f52d70",
  1739 => x"84808029",
  1740 => x"1280def3",
  1741 => x"0b80f52d",
  1742 => x"70982b81",
  1743 => x"f00a0672",
  1744 => x"057080e6",
  1745 => x"e40cfe11",
  1746 => x"7e297705",
  1747 => x"80e6e80c",
  1748 => x"52595243",
  1749 => x"545e5152",
  1750 => x"59525d57",
  1751 => x"5957b7b9",
  1752 => x"0480ded6",
  1753 => x"0b80f52d",
  1754 => x"80ded50b",
  1755 => x"80f52d71",
  1756 => x"82802905",
  1757 => x"7080e6d8",
  1758 => x"0c70a029",
  1759 => x"83ff0570",
  1760 => x"892a7080",
  1761 => x"e6ec0c80",
  1762 => x"dedb0b80",
  1763 => x"f52d80de",
  1764 => x"da0b80f5",
  1765 => x"2d718280",
  1766 => x"29057080",
  1767 => x"e6f40c7b",
  1768 => x"71291e70",
  1769 => x"80e6e80c",
  1770 => x"7d80e6e4",
  1771 => x"0c730580",
  1772 => x"e6e00c55",
  1773 => x"5e515155",
  1774 => x"558051b0",
  1775 => x"902d8155",
  1776 => x"7480ddcc",
  1777 => x"0c02a805",
  1778 => x"0d0402ec",
  1779 => x"050d7670",
  1780 => x"872c7180",
  1781 => x"ff065556",
  1782 => x"5480e6d4",
  1783 => x"088a3873",
  1784 => x"882c7481",
  1785 => x"ff065455",
  1786 => x"80dec452",
  1787 => x"80e6dc08",
  1788 => x"1551aead",
  1789 => x"2d80ddcc",
  1790 => x"085480dd",
  1791 => x"cc08802e",
  1792 => x"b83880e6",
  1793 => x"d408802e",
  1794 => x"9a387284",
  1795 => x"2980dec4",
  1796 => x"05700852",
  1797 => x"53beb12d",
  1798 => x"80ddcc08",
  1799 => x"f00a0653",
  1800 => x"b8b70472",
  1801 => x"1080dec4",
  1802 => x"057080e0",
  1803 => x"2d5253be",
  1804 => x"e22d80dd",
  1805 => x"cc085372",
  1806 => x"547380dd",
  1807 => x"cc0c0294",
  1808 => x"050d0402",
  1809 => x"e4050d78",
  1810 => x"70842c80",
  1811 => x"e6fc0805",
  1812 => x"718f0652",
  1813 => x"5553728a",
  1814 => x"3880dec4",
  1815 => x"527351ae",
  1816 => x"ad2d72a0",
  1817 => x"2980dec4",
  1818 => x"05558075",
  1819 => x"80f52d57",
  1820 => x"5375732e",
  1821 => x"83388153",
  1822 => x"7581e52e",
  1823 => x"828b3881",
  1824 => x"70740654",
  1825 => x"5772802e",
  1826 => x"81ff388b",
  1827 => x"1580f52d",
  1828 => x"70832a70",
  1829 => x"79065154",
  1830 => x"54729b38",
  1831 => x"80dc9008",
  1832 => x"54738938",
  1833 => x"7380e2c4",
  1834 => x"0b81b72d",
  1835 => x"7280dc90",
  1836 => x"0c7453bb",
  1837 => x"8b04738f",
  1838 => x"2e098106",
  1839 => x"81cb3875",
  1840 => x"9f068d29",
  1841 => x"80e2b705",
  1842 => x"54811580",
  1843 => x"f52d7470",
  1844 => x"81055681",
  1845 => x"b72d8315",
  1846 => x"80f52d74",
  1847 => x"70810556",
  1848 => x"81b72d85",
  1849 => x"1580f52d",
  1850 => x"74708105",
  1851 => x"5681b72d",
  1852 => x"871580f5",
  1853 => x"2d747081",
  1854 => x"055681b7",
  1855 => x"2d891580",
  1856 => x"f52d7470",
  1857 => x"81055681",
  1858 => x"b72d8e15",
  1859 => x"80f52d74",
  1860 => x"70810556",
  1861 => x"81b72d90",
  1862 => x"1580f52d",
  1863 => x"74708105",
  1864 => x"5681b72d",
  1865 => x"921580f5",
  1866 => x"2d747081",
  1867 => x"055681b7",
  1868 => x"2d941580",
  1869 => x"f52d7470",
  1870 => x"81055681",
  1871 => x"b72d9615",
  1872 => x"80f52d74",
  1873 => x"70810556",
  1874 => x"81b72d98",
  1875 => x"1580f52d",
  1876 => x"74708105",
  1877 => x"5681b72d",
  1878 => x"9c1580f5",
  1879 => x"2d747081",
  1880 => x"055681b7",
  1881 => x"2d9e1580",
  1882 => x"f52d7470",
  1883 => x"81055681",
  1884 => x"b72d7586",
  1885 => x"2a708106",
  1886 => x"51537280",
  1887 => x"2e863880",
  1888 => x"7481b72d",
  1889 => x"7680dc90",
  1890 => x"0c805372",
  1891 => x"80ddcc0c",
  1892 => x"029c050d",
  1893 => x"0402cc05",
  1894 => x"0d7e605e",
  1895 => x"5b800b80",
  1896 => x"e6f80880",
  1897 => x"e6fc0859",
  1898 => x"5d568059",
  1899 => x"80e6d808",
  1900 => x"792e81de",
  1901 => x"38788f06",
  1902 => x"a0175754",
  1903 => x"73913880",
  1904 => x"dec45276",
  1905 => x"51811757",
  1906 => x"aead2d80",
  1907 => x"dec45680",
  1908 => x"7680f52d",
  1909 => x"56547474",
  1910 => x"2e833881",
  1911 => x"547481e5",
  1912 => x"2e81a338",
  1913 => x"81707506",
  1914 => x"555a7380",
  1915 => x"2e819738",
  1916 => x"8b1680f5",
  1917 => x"2d709806",
  1918 => x"59547780",
  1919 => x"e3388b53",
  1920 => x"7c527551",
  1921 => x"afd12d80",
  1922 => x"ddcc0880",
  1923 => x"f9389c16",
  1924 => x"0851beb1",
  1925 => x"2d80ddcc",
  1926 => x"08841c0c",
  1927 => x"9a1680e0",
  1928 => x"2d51bee2",
  1929 => x"2d80ddcc",
  1930 => x"0880ddcc",
  1931 => x"08881d0c",
  1932 => x"80ddcc08",
  1933 => x"555580e6",
  1934 => x"d408802e",
  1935 => x"99389416",
  1936 => x"80e02d51",
  1937 => x"bee22d80",
  1938 => x"ddcc0890",
  1939 => x"2b83fff0",
  1940 => x"0a067016",
  1941 => x"51547388",
  1942 => x"1c0c777b",
  1943 => x"0cbd8104",
  1944 => x"73842a70",
  1945 => x"81065154",
  1946 => x"73802e9a",
  1947 => x"388b537c",
  1948 => x"527551af",
  1949 => x"d12d80dd",
  1950 => x"cc088b38",
  1951 => x"7551b090",
  1952 => x"2d7954bd",
  1953 => x"ce048119",
  1954 => x"5980e6d8",
  1955 => x"087926fe",
  1956 => x"a43880e6",
  1957 => x"d408802e",
  1958 => x"b3387b51",
  1959 => x"b7ca2d80",
  1960 => x"ddcc0880",
  1961 => x"ddcc0880",
  1962 => x"fffffff8",
  1963 => x"06555c73",
  1964 => x"80ffffff",
  1965 => x"f82e9538",
  1966 => x"80ddcc08",
  1967 => x"fe0580e6",
  1968 => x"cc082980",
  1969 => x"e6e00805",
  1970 => x"57bbaa04",
  1971 => x"80547380",
  1972 => x"ddcc0c02",
  1973 => x"b4050d04",
  1974 => x"02f4050d",
  1975 => x"74700881",
  1976 => x"05710c70",
  1977 => x"0880e6d0",
  1978 => x"08065353",
  1979 => x"718f3888",
  1980 => x"130851b7",
  1981 => x"ca2d80dd",
  1982 => x"cc088814",
  1983 => x"0c810b80",
  1984 => x"ddcc0c02",
  1985 => x"8c050d04",
  1986 => x"02f0050d",
  1987 => x"75881108",
  1988 => x"fe0580e6",
  1989 => x"cc082980",
  1990 => x"e6e00811",
  1991 => x"720880e6",
  1992 => x"d0080605",
  1993 => x"79555354",
  1994 => x"54aead2d",
  1995 => x"0290050d",
  1996 => x"0402f405",
  1997 => x"0d747088",
  1998 => x"2a83fe80",
  1999 => x"06707298",
  2000 => x"2a077288",
  2001 => x"2b87fc80",
  2002 => x"80067398",
  2003 => x"2b81f00a",
  2004 => x"06717307",
  2005 => x"0780ddcc",
  2006 => x"0c565153",
  2007 => x"51028c05",
  2008 => x"0d0402f8",
  2009 => x"050d028e",
  2010 => x"0580f52d",
  2011 => x"74882b07",
  2012 => x"7083ffff",
  2013 => x"0680ddcc",
  2014 => x"0c510288",
  2015 => x"050d0402",
  2016 => x"ec050d76",
  2017 => x"787a5355",
  2018 => x"52815580",
  2019 => x"7125ae38",
  2020 => x"70537370",
  2021 => x"81055580",
  2022 => x"f52d7270",
  2023 => x"81055481",
  2024 => x"b72d7380",
  2025 => x"f52d5170",
  2026 => x"86387055",
  2027 => x"bfb20474",
  2028 => x"8638a072",
  2029 => x"81b72dff",
  2030 => x"135372d6",
  2031 => x"38807270",
  2032 => x"81055481",
  2033 => x"b72d8072",
  2034 => x"81b72d02",
  2035 => x"94050d04",
  2036 => x"02e8050d",
  2037 => x"77568070",
  2038 => x"56547376",
  2039 => x"24b63880",
  2040 => x"e6d80874",
  2041 => x"2eae3873",
  2042 => x"51b8c32d",
  2043 => x"80ddcc08",
  2044 => x"80ddcc08",
  2045 => x"09810570",
  2046 => x"80ddcc08",
  2047 => x"079f2a77",
  2048 => x"05811757",
  2049 => x"57535374",
  2050 => x"76248938",
  2051 => x"80e6d808",
  2052 => x"7426d438",
  2053 => x"7280ddcc",
  2054 => x"0c029805",
  2055 => x"0d0402f0",
  2056 => x"050d80dd",
  2057 => x"c8081651",
  2058 => x"bfd02d80",
  2059 => x"ddcc0854",
  2060 => x"80ddcc08",
  2061 => x"802ebb38",
  2062 => x"8b5380dd",
  2063 => x"cc085280",
  2064 => x"e2c451be",
  2065 => x"ff2d8853",
  2066 => x"735280e4",
  2067 => x"c851beff",
  2068 => x"2d835380",
  2069 => x"d3cc5280",
  2070 => x"e4d051be",
  2071 => x"ff2d80e7",
  2072 => x"84085473",
  2073 => x"802e8b38",
  2074 => x"80e4c852",
  2075 => x"80e2c451",
  2076 => x"732d0290",
  2077 => x"050d0402",
  2078 => x"dc050d80",
  2079 => x"705a5574",
  2080 => x"80ddc808",
  2081 => x"25b43880",
  2082 => x"e6d80875",
  2083 => x"2eac3878",
  2084 => x"51b8c32d",
  2085 => x"80ddcc08",
  2086 => x"09810570",
  2087 => x"80ddcc08",
  2088 => x"079f2a76",
  2089 => x"05811b5b",
  2090 => x"56547480",
  2091 => x"ddc80825",
  2092 => x"893880e6",
  2093 => x"d8087926",
  2094 => x"d6388055",
  2095 => x"7880e6d8",
  2096 => x"082781e2",
  2097 => x"387851b8",
  2098 => x"c32d80dd",
  2099 => x"cc08802e",
  2100 => x"81b33880",
  2101 => x"ddcc088b",
  2102 => x"0580f52d",
  2103 => x"70842a70",
  2104 => x"81067710",
  2105 => x"78842b80",
  2106 => x"e2c40b80",
  2107 => x"f52d5c5c",
  2108 => x"53515556",
  2109 => x"73802e80",
  2110 => x"ce387416",
  2111 => x"822b80c3",
  2112 => x"ca0b80dc",
  2113 => x"9c120c54",
  2114 => x"77753110",
  2115 => x"80e78811",
  2116 => x"55569074",
  2117 => x"70810556",
  2118 => x"81b72da0",
  2119 => x"7481b72d",
  2120 => x"7681ff06",
  2121 => x"81165854",
  2122 => x"73802e8b",
  2123 => x"389c5380",
  2124 => x"e2c45280",
  2125 => x"c2be048b",
  2126 => x"5380ddcc",
  2127 => x"085280e7",
  2128 => x"8a165180",
  2129 => x"c2fc0474",
  2130 => x"16822b80",
  2131 => x"c09e0b80",
  2132 => x"dc9c120c",
  2133 => x"547681ff",
  2134 => x"06811658",
  2135 => x"5473802e",
  2136 => x"8b389c53",
  2137 => x"80e2c452",
  2138 => x"80c2f304",
  2139 => x"8b5380dd",
  2140 => x"cc085277",
  2141 => x"75311080",
  2142 => x"e7880551",
  2143 => x"7655beff",
  2144 => x"2d80c39a",
  2145 => x"04749029",
  2146 => x"75317010",
  2147 => x"80e78805",
  2148 => x"515480dd",
  2149 => x"cc087481",
  2150 => x"b72d8119",
  2151 => x"59748b24",
  2152 => x"a43880c1",
  2153 => x"bc047490",
  2154 => x"29753170",
  2155 => x"1080e788",
  2156 => x"058c7731",
  2157 => x"57515480",
  2158 => x"7481b72d",
  2159 => x"9e14ff16",
  2160 => x"565474f3",
  2161 => x"3802a405",
  2162 => x"0d0402fc",
  2163 => x"050d80dd",
  2164 => x"c8081351",
  2165 => x"bfd02d80",
  2166 => x"ddcc0880",
  2167 => x"2e893880",
  2168 => x"ddcc0851",
  2169 => x"b0902d80",
  2170 => x"0b80ddc8",
  2171 => x"0c80c0f7",
  2172 => x"2d99ed2d",
  2173 => x"0284050d",
  2174 => x"0402f805",
  2175 => x"0d735170",
  2176 => x"fd2eb338",
  2177 => x"70fd248b",
  2178 => x"3870fc2e",
  2179 => x"80d13880",
  2180 => x"c4f90470",
  2181 => x"fe2eba38",
  2182 => x"70ff2e09",
  2183 => x"810680d9",
  2184 => x"3880ddc8",
  2185 => x"08517080",
  2186 => x"2e80ce38",
  2187 => x"ff1180dd",
  2188 => x"c80c80c4",
  2189 => x"f90480dd",
  2190 => x"c808f405",
  2191 => x"7080ddc8",
  2192 => x"0c517080",
  2193 => x"25b33880",
  2194 => x"0b80ddc8",
  2195 => x"0c80c4f9",
  2196 => x"0480ddc8",
  2197 => x"08810580",
  2198 => x"ddc80c80",
  2199 => x"c4f90480",
  2200 => x"ddc8088c",
  2201 => x"117080dd",
  2202 => x"c80c5252",
  2203 => x"80e6d808",
  2204 => x"71268638",
  2205 => x"7180ddc8",
  2206 => x"0c80c0f7",
  2207 => x"2d99ed2d",
  2208 => x"0288050d",
  2209 => x"0402fc05",
  2210 => x"0d800b80",
  2211 => x"ddc80c80",
  2212 => x"c0f72d98",
  2213 => x"d62d80dd",
  2214 => x"cc0880dd",
  2215 => x"b80c80dc",
  2216 => x"94519b93",
  2217 => x"2d028405",
  2218 => x"0d0402f8",
  2219 => x"050d810b",
  2220 => x"80d5dc0c",
  2221 => x"80ddf408",
  2222 => x"bff9ff06",
  2223 => x"81800770",
  2224 => x"80ddf40c",
  2225 => x"fc0c7351",
  2226 => x"80c5852d",
  2227 => x"0288050d",
  2228 => x"0402f805",
  2229 => x"0d820b80",
  2230 => x"d5dc0c80",
  2231 => x"ddf408bf",
  2232 => x"faff0682",
  2233 => x"80077080",
  2234 => x"ddf40cfc",
  2235 => x"0c735180",
  2236 => x"c5852d02",
  2237 => x"88050d04",
  2238 => x"02f8050d",
  2239 => x"830b80d5",
  2240 => x"dc0c80dd",
  2241 => x"f408bfff",
  2242 => x"ff068780",
  2243 => x"077080dd",
  2244 => x"f40cfc0c",
  2245 => x"735180c5",
  2246 => x"852d0288",
  2247 => x"050d0471",
  2248 => x"80e7840c",
  2249 => x"04000000",
  2250 => x"00ffffff",
  2251 => x"ff00ffff",
  2252 => x"ffff00ff",
  2253 => x"ffffff00",
  2254 => x"434f4e46",
  2255 => x"49472020",
  2256 => x"54585400",
  2257 => x"00000000",
  2258 => x"54686572",
  2259 => x"65206973",
  2260 => x"206e6f20",
  2261 => x"696d6167",
  2262 => x"65207768",
  2263 => x"656e206c",
  2264 => x"6f616469",
  2265 => x"6e670000",
  2266 => x"436f6e74",
  2267 => x"696e7565",
  2268 => x"00000000",
  2269 => x"3d205a58",
  2270 => x"38312f5a",
  2271 => x"58383020",
  2272 => x"436f6e66",
  2273 => x"69677572",
  2274 => x"6174696f",
  2275 => x"6e203d00",
  2276 => x"3d3d3d3d",
  2277 => x"3d3d3d3d",
  2278 => x"3d3d3d3d",
  2279 => x"3d3d3d3d",
  2280 => x"3d3d3d3d",
  2281 => x"3d3d3d3d",
  2282 => x"3d3d3d00",
  2283 => x"4c6f7720",
  2284 => x"52414d3a",
  2285 => x"204f6666",
  2286 => x"2f384b42",
  2287 => x"00000000",
  2288 => x"51532043",
  2289 => x"4852533a",
  2290 => x"44697361",
  2291 => x"626c6564",
  2292 => x"2f456e61",
  2293 => x"626c6564",
  2294 => x"28463129",
  2295 => x"00000000",
  2296 => x"4348524f",
  2297 => x"4d413831",
  2298 => x"3a204469",
  2299 => x"7361626c",
  2300 => x"65642f45",
  2301 => x"6e61626c",
  2302 => x"65640000",
  2303 => x"496e7665",
  2304 => x"72736520",
  2305 => x"76696465",
  2306 => x"6f3a204f",
  2307 => x"66662f4f",
  2308 => x"6e000000",
  2309 => x"426c6163",
  2310 => x"6b20626f",
  2311 => x"72646572",
  2312 => x"3a204f66",
  2313 => x"662f4f6e",
  2314 => x"00000000",
  2315 => x"56696465",
  2316 => x"6f206672",
  2317 => x"65717565",
  2318 => x"6e63793a",
  2319 => x"20353048",
  2320 => x"7a2f3630",
  2321 => x"487a0000",
  2322 => x"476f2042",
  2323 => x"61636b00",
  2324 => x"536c6f77",
  2325 => x"206d6f64",
  2326 => x"65207370",
  2327 => x"6565643a",
  2328 => x"204f7269",
  2329 => x"67696e61",
  2330 => x"6c000000",
  2331 => x"536c6f77",
  2332 => x"206d6f64",
  2333 => x"65207370",
  2334 => x"6565643a",
  2335 => x"204e6f57",
  2336 => x"61697400",
  2337 => x"536c6f77",
  2338 => x"206d6f64",
  2339 => x"65207370",
  2340 => x"6565643a",
  2341 => x"20783200",
  2342 => x"536c6f77",
  2343 => x"206d6f64",
  2344 => x"65207370",
  2345 => x"6565643a",
  2346 => x"20783800",
  2347 => x"43485224",
  2348 => x"3132382f",
  2349 => x"5544473a",
  2350 => x"20313238",
  2351 => x"20436861",
  2352 => x"72730000",
  2353 => x"43485224",
  2354 => x"3132382f",
  2355 => x"5544473a",
  2356 => x"20363420",
  2357 => x"43686172",
  2358 => x"73000000",
  2359 => x"43485224",
  2360 => x"3132382f",
  2361 => x"5544473a",
  2362 => x"20446973",
  2363 => x"61626c65",
  2364 => x"64000000",
  2365 => x"4a6f7973",
  2366 => x"7469636b",
  2367 => x"3a204375",
  2368 => x"72736f72",
  2369 => x"00000000",
  2370 => x"4a6f7973",
  2371 => x"7469636b",
  2372 => x"3a205369",
  2373 => x"6e636c61",
  2374 => x"69720000",
  2375 => x"4a6f7973",
  2376 => x"7469636b",
  2377 => x"3a205a58",
  2378 => x"38310000",
  2379 => x"4d61696e",
  2380 => x"2052414d",
  2381 => x"3a203136",
  2382 => x"4b420000",
  2383 => x"4d61696e",
  2384 => x"2052414d",
  2385 => x"3a203332",
  2386 => x"4b420000",
  2387 => x"4d61696e",
  2388 => x"2052414d",
  2389 => x"3a203438",
  2390 => x"4b420000",
  2391 => x"4d61696e",
  2392 => x"2052414d",
  2393 => x"3a20314b",
  2394 => x"42000000",
  2395 => x"436f6d70",
  2396 => x"75746572",
  2397 => x"204d6f64",
  2398 => x"656c3a20",
  2399 => x"5a583831",
  2400 => x"00000000",
  2401 => x"436f6d70",
  2402 => x"75746572",
  2403 => x"204d6f64",
  2404 => x"656c3a20",
  2405 => x"5a583830",
  2406 => x"00000000",
  2407 => x"3d3d205a",
  2408 => x"5838312f",
  2409 => x"5a583830",
  2410 => x"20666f72",
  2411 => x"205a5844",
  2412 => x"4f53203d",
  2413 => x"3d000000",
  2414 => x"3d3d3d3d",
  2415 => x"3d3d3d3d",
  2416 => x"3d3d3d3d",
  2417 => x"3d3d3d3d",
  2418 => x"3d3d3d3d",
  2419 => x"3d3d3d3d",
  2420 => x"3d000000",
  2421 => x"52657365",
  2422 => x"74000000",
  2423 => x"4c6f6164",
  2424 => x"20546170",
  2425 => x"6520282e",
  2426 => x"70292010",
  2427 => x"00000000",
  2428 => x"4c6f6164",
  2429 => x"20546170",
  2430 => x"6520282e",
  2431 => x"6f292010",
  2432 => x"00000000",
  2433 => x"4c6f6164",
  2434 => x"20526f6d",
  2435 => x"2020282e",
  2436 => x"726f6d29",
  2437 => x"20100000",
  2438 => x"436f6e66",
  2439 => x"69677572",
  2440 => x"6174696f",
  2441 => x"6e206f70",
  2442 => x"74696f6e",
  2443 => x"73201000",
  2444 => x"4b657962",
  2445 => x"6f617264",
  2446 => x"2048656c",
  2447 => x"70000000",
  2448 => x"45786974",
  2449 => x"00000000",
  2450 => x"3d3d205a",
  2451 => x"5838312f",
  2452 => x"5a583830",
  2453 => x"20666f72",
  2454 => x"205a5855",
  2455 => x"4e4f203d",
  2456 => x"3d000000",
  2457 => x"524f4d20",
  2458 => x"6c6f6164",
  2459 => x"696e6720",
  2460 => x"6661696c",
  2461 => x"65640000",
  2462 => x"4f4b0000",
  2463 => x"54617065",
  2464 => x"2066696c",
  2465 => x"65204c6f",
  2466 => x"61646564",
  2467 => x"2e000000",
  2468 => x"54797065",
  2469 => x"204c4f41",
  2470 => x"44202222",
  2471 => x"202b2045",
  2472 => x"4e544552",
  2473 => x"206f6e20",
  2474 => x"5a583831",
  2475 => x"00000000",
  2476 => x"3d205a58",
  2477 => x"38312f5a",
  2478 => x"58383020",
  2479 => x"4b657962",
  2480 => x"6f617264",
  2481 => x"2048656c",
  2482 => x"70203d00",
  2483 => x"5363726f",
  2484 => x"6c6c204c",
  2485 => x"6f636b3a",
  2486 => x"20636861",
  2487 => x"6e676520",
  2488 => x"62657477",
  2489 => x"65656e00",
  2490 => x"52474220",
  2491 => x"616e6420",
  2492 => x"56474120",
  2493 => x"76696465",
  2494 => x"6f206d6f",
  2495 => x"64650000",
  2496 => x"4374726c",
  2497 => x"2b416c74",
  2498 => x"2b44656c",
  2499 => x"6574653a",
  2500 => x"20536f66",
  2501 => x"74205265",
  2502 => x"73657400",
  2503 => x"4374726c",
  2504 => x"2b416c74",
  2505 => x"2b426163",
  2506 => x"6b737061",
  2507 => x"63653a20",
  2508 => x"48617264",
  2509 => x"20726573",
  2510 => x"65740000",
  2511 => x"4635206f",
  2512 => x"72206a6f",
  2513 => x"79737469",
  2514 => x"636b2062",
  2515 => x"742e323a",
  2516 => x"20746f20",
  2517 => x"73686f77",
  2518 => x"00000000",
  2519 => x"6f722068",
  2520 => x"69646520",
  2521 => x"74686520",
  2522 => x"6f707469",
  2523 => x"6f6e7320",
  2524 => x"6d656e75",
  2525 => x"2e000000",
  2526 => x"57415344",
  2527 => x"202f2063",
  2528 => x"7572736f",
  2529 => x"72206b65",
  2530 => x"7973202f",
  2531 => x"206a6f79",
  2532 => x"73746963",
  2533 => x"6b000000",
  2534 => x"746f2073",
  2535 => x"656c6563",
  2536 => x"74206d65",
  2537 => x"6e75206f",
  2538 => x"7074696f",
  2539 => x"6e2e0000",
  2540 => x"456e7465",
  2541 => x"72202f20",
  2542 => x"46697265",
  2543 => x"20746f20",
  2544 => x"63686f6f",
  2545 => x"7365206f",
  2546 => x"7074696f",
  2547 => x"6e2e0000",
  2548 => x"3d205a58",
  2549 => x"38312f5a",
  2550 => x"58383020",
  2551 => x"436f7265",
  2552 => x"20437265",
  2553 => x"64697473",
  2554 => x"20203d00",
  2555 => x"5a583831",
  2556 => x"2f5a5838",
  2557 => x"3020636f",
  2558 => x"72652066",
  2559 => x"6f72205a",
  2560 => x"58554e4f",
  2561 => x"2c200000",
  2562 => x"5a58444f",
  2563 => x"5320616e",
  2564 => x"64205a58",
  2565 => x"444f532b",
  2566 => x"20626f61",
  2567 => x"7264732e",
  2568 => x"00000000",
  2569 => x"4f726967",
  2570 => x"696e616c",
  2571 => x"20636f72",
  2572 => x"65732062",
  2573 => x"793a0000",
  2574 => x"202d2053",
  2575 => x"7a6f6d62",
  2576 => x"61746865",
  2577 => x"6c796920",
  2578 => x"47796f72",
  2579 => x"67792028",
  2580 => x"4d697374",
  2581 => x"29000000",
  2582 => x"202d2053",
  2583 => x"6f726765",
  2584 => x"6c696720",
  2585 => x"284d6973",
  2586 => x"74657229",
  2587 => x"00000000",
  2588 => x"202d204a",
  2589 => x"6f746567",
  2590 => x"6f20284a",
  2591 => x"54343920",
  2592 => x"64656769",
  2593 => x"676e2900",
  2594 => x"506f7274",
  2595 => x"206d6164",
  2596 => x"65206279",
  2597 => x"3a204176",
  2598 => x"6c697841",
  2599 => x"00000000",
  2600 => x"496e6974",
  2601 => x"69616c69",
  2602 => x"7a696e67",
  2603 => x"20534420",
  2604 => x"63617264",
  2605 => x"0a000000",
  2606 => x"4c6f6164",
  2607 => x"696e6720",
  2608 => x"696e6974",
  2609 => x"69616c20",
  2610 => x"524f4d2e",
  2611 => x"2e2e0a00",
  2612 => x"5a583831",
  2613 => x"20202020",
  2614 => x"20202000",
  2615 => x"524f4d53",
  2616 => x"20202020",
  2617 => x"20202000",
  2618 => x"5a583858",
  2619 => x"20202020",
  2620 => x"524f4d00",
  2621 => x"4572726f",
  2622 => x"72204c6f",
  2623 => x"6164696e",
  2624 => x"6720524f",
  2625 => x"4d2e2e2e",
  2626 => x"0a000000",
  2627 => x"2e2e2020",
  2628 => x"20202020",
  2629 => x"20202000",
  2630 => x"16200000",
  2631 => x"14200000",
  2632 => x"15200000",
  2633 => x"53442069",
  2634 => x"6e69742e",
  2635 => x"2e2e0a00",
  2636 => x"53442063",
  2637 => x"61726420",
  2638 => x"72657365",
  2639 => x"74206661",
  2640 => x"696c6564",
  2641 => x"210a0000",
  2642 => x"53444843",
  2643 => x"20657272",
  2644 => x"6f72210a",
  2645 => x"00000000",
  2646 => x"57726974",
  2647 => x"65206661",
  2648 => x"696c6564",
  2649 => x"0a000000",
  2650 => x"52656164",
  2651 => x"20666169",
  2652 => x"6c65640a",
  2653 => x"00000000",
  2654 => x"43617264",
  2655 => x"20696e69",
  2656 => x"74206661",
  2657 => x"696c6564",
  2658 => x"0a000000",
  2659 => x"46415431",
  2660 => x"36202020",
  2661 => x"00000000",
  2662 => x"46415433",
  2663 => x"32202020",
  2664 => x"00000000",
  2665 => x"4e6f2070",
  2666 => x"61727469",
  2667 => x"74696f6e",
  2668 => x"20736967",
  2669 => x"0a000000",
  2670 => x"42616420",
  2671 => x"70617274",
  2672 => x"0a000000",
  2673 => x"4261636b",
  2674 => x"00000000",
  2675 => x"434f4c00",
  2676 => x"00000002",
  2677 => x"00000002",
  2678 => x"00002374",
  2679 => x"00000342",
  2680 => x"00000002",
  2681 => x"00002390",
  2682 => x"00000342",
  2683 => x"00000003",
  2684 => x"00002ac0",
  2685 => x"00000002",
  2686 => x"00000003",
  2687 => x"00002ab0",
  2688 => x"00000004",
  2689 => x"00000001",
  2690 => x"000023ac",
  2691 => x"00000000",
  2692 => x"00000003",
  2693 => x"00002aa4",
  2694 => x"00000003",
  2695 => x"00000001",
  2696 => x"000023c0",
  2697 => x"00000001",
  2698 => x"00000003",
  2699 => x"00002a98",
  2700 => x"00000003",
  2701 => x"00000001",
  2702 => x"000023e0",
  2703 => x"00000002",
  2704 => x"00000001",
  2705 => x"000023fc",
  2706 => x"00000003",
  2707 => x"00000001",
  2708 => x"00002414",
  2709 => x"00000004",
  2710 => x"00000003",
  2711 => x"00002a88",
  2712 => x"00000003",
  2713 => x"00000001",
  2714 => x"0000242c",
  2715 => x"00000005",
  2716 => x"00000004",
  2717 => x"00002448",
  2718 => x"00002ef8",
  2719 => x"00000000",
  2720 => x"00000000",
  2721 => x"00000000",
  2722 => x"00002450",
  2723 => x"0000246c",
  2724 => x"00002484",
  2725 => x"00002498",
  2726 => x"000024ac",
  2727 => x"000024c4",
  2728 => x"000024dc",
  2729 => x"000024f4",
  2730 => x"00002508",
  2731 => x"0000251c",
  2732 => x"0000252c",
  2733 => x"0000253c",
  2734 => x"0000254c",
  2735 => x"0000255c",
  2736 => x"0000256c",
  2737 => x"00002584",
  2738 => x"30303030",
  2739 => x"30303030",
  2740 => x"30303030",
  2741 => x"00000000",
  2742 => x"00000000",
  2743 => x"00000000",
  2744 => x"00000002",
  2745 => x"0000259c",
  2746 => x"00000343",
  2747 => x"00000002",
  2748 => x"000025b8",
  2749 => x"00000343",
  2750 => x"00000002",
  2751 => x"000025d4",
  2752 => x"00000386",
  2753 => x"00000002",
  2754 => x"000025dc",
  2755 => x"000022aa",
  2756 => x"00000002",
  2757 => x"000025f0",
  2758 => x"000022d1",
  2759 => x"00000002",
  2760 => x"00002604",
  2761 => x"000022f8",
  2762 => x"00000002",
  2763 => x"00002618",
  2764 => x"00000353",
  2765 => x"00000002",
  2766 => x"00002630",
  2767 => x"00000363",
  2768 => x"00000002",
  2769 => x"00002640",
  2770 => x"00000c73",
  2771 => x"00000000",
  2772 => x"00000000",
  2773 => x"00000000",
  2774 => x"00000002",
  2775 => x"00002648",
  2776 => x"00000343",
  2777 => x"00000002",
  2778 => x"000025b8",
  2779 => x"00000343",
  2780 => x"00000002",
  2781 => x"000025d4",
  2782 => x"00000386",
  2783 => x"00000002",
  2784 => x"000025dc",
  2785 => x"000022aa",
  2786 => x"00000002",
  2787 => x"000025f0",
  2788 => x"000022d1",
  2789 => x"00000002",
  2790 => x"00002604",
  2791 => x"000022f8",
  2792 => x"00000002",
  2793 => x"00002618",
  2794 => x"00000353",
  2795 => x"00000002",
  2796 => x"00002630",
  2797 => x"00000363",
  2798 => x"00000002",
  2799 => x"00002640",
  2800 => x"00000c73",
  2801 => x"00000000",
  2802 => x"00000000",
  2803 => x"00000000",
  2804 => x"00000004",
  2805 => x"00002664",
  2806 => x"00002bd0",
  2807 => x"00000004",
  2808 => x"00002678",
  2809 => x"00002ef8",
  2810 => x"00000000",
  2811 => x"00000000",
  2812 => x"00000000",
  2813 => x"00000004",
  2814 => x"0000267c",
  2815 => x"00002bf4",
  2816 => x"00000004",
  2817 => x"00002690",
  2818 => x"00002bf4",
  2819 => x"00000004",
  2820 => x"00002954",
  2821 => x"00002bf4",
  2822 => x"00000004",
  2823 => x"00002348",
  2824 => x"00002bf4",
  2825 => x"00000004",
  2826 => x"00002954",
  2827 => x"00002bf4",
  2828 => x"00000004",
  2829 => x"00002368",
  2830 => x"00002ef8",
  2831 => x"00000000",
  2832 => x"00000000",
  2833 => x"00000000",
  2834 => x"00000002",
  2835 => x"000026b0",
  2836 => x"00000342",
  2837 => x"00000002",
  2838 => x"00002390",
  2839 => x"00000342",
  2840 => x"00000002",
  2841 => x"000026cc",
  2842 => x"00000342",
  2843 => x"00000002",
  2844 => x"000026e8",
  2845 => x"00000342",
  2846 => x"00000002",
  2847 => x"00002700",
  2848 => x"00000342",
  2849 => x"00000002",
  2850 => x"0000271c",
  2851 => x"00000342",
  2852 => x"00000002",
  2853 => x"0000273c",
  2854 => x"00000342",
  2855 => x"00000002",
  2856 => x"0000275c",
  2857 => x"00000342",
  2858 => x"00000002",
  2859 => x"00002778",
  2860 => x"00000342",
  2861 => x"00000002",
  2862 => x"00002798",
  2863 => x"00000342",
  2864 => x"00000002",
  2865 => x"000027b0",
  2866 => x"00000342",
  2867 => x"00000002",
  2868 => x"00002954",
  2869 => x"00000342",
  2870 => x"00000004",
  2871 => x"00002678",
  2872 => x"00002ef8",
  2873 => x"00000000",
  2874 => x"00000000",
  2875 => x"00000000",
  2876 => x"00000002",
  2877 => x"000027d0",
  2878 => x"00000342",
  2879 => x"00000002",
  2880 => x"00002390",
  2881 => x"00000342",
  2882 => x"00000002",
  2883 => x"000027ec",
  2884 => x"00000342",
  2885 => x"00000002",
  2886 => x"00002808",
  2887 => x"00000342",
  2888 => x"00000002",
  2889 => x"00002954",
  2890 => x"00000342",
  2891 => x"00000002",
  2892 => x"00002824",
  2893 => x"00000342",
  2894 => x"00000002",
  2895 => x"00002838",
  2896 => x"00000342",
  2897 => x"00000002",
  2898 => x"00002858",
  2899 => x"00000342",
  2900 => x"00000002",
  2901 => x"00002870",
  2902 => x"00000342",
  2903 => x"00000002",
  2904 => x"00002954",
  2905 => x"00000342",
  2906 => x"00000002",
  2907 => x"00002888",
  2908 => x"00000342",
  2909 => x"00000002",
  2910 => x"00002954",
  2911 => x"00000342",
  2912 => x"00000004",
  2913 => x"00002678",
  2914 => x"00002ef8",
  2915 => x"00000000",
  2916 => x"00000000",
  2917 => x"00000000",
  2918 => x"00000000",
  2919 => x"00000000",
  2920 => x"00000000",
  2921 => x"00000000",
  2922 => x"00000000",
  2923 => x"00000000",
  2924 => x"00000000",
  2925 => x"00000000",
  2926 => x"00000000",
  2927 => x"00000000",
  2928 => x"00000000",
  2929 => x"00000000",
  2930 => x"00000000",
  2931 => x"00000000",
  2932 => x"00000000",
  2933 => x"00000000",
  2934 => x"00000000",
  2935 => x"00000000",
  2936 => x"00000006",
  2937 => x"00000043",
  2938 => x"00000042",
  2939 => x"0000003b",
  2940 => x"0000004b",
  2941 => x"0000007e",
  2942 => x"00000003",
  2943 => x"0000000b",
  2944 => x"00000083",
  2945 => x"00000023",
  2946 => x"0000007e",
  2947 => x"00000000",
  2948 => x"00000000",
  2949 => x"00000002",
  2950 => x"00003388",
  2951 => x"0000201e",
  2952 => x"00000002",
  2953 => x"000033a6",
  2954 => x"0000201e",
  2955 => x"00000002",
  2956 => x"000033c4",
  2957 => x"0000201e",
  2958 => x"00000002",
  2959 => x"000033e2",
  2960 => x"0000201e",
  2961 => x"00000002",
  2962 => x"00003400",
  2963 => x"0000201e",
  2964 => x"00000002",
  2965 => x"0000341e",
  2966 => x"0000201e",
  2967 => x"00000002",
  2968 => x"0000343c",
  2969 => x"0000201e",
  2970 => x"00000002",
  2971 => x"0000345a",
  2972 => x"0000201e",
  2973 => x"00000002",
  2974 => x"00003478",
  2975 => x"0000201e",
  2976 => x"00000002",
  2977 => x"00003496",
  2978 => x"0000201e",
  2979 => x"00000002",
  2980 => x"000034b4",
  2981 => x"0000201e",
  2982 => x"00000002",
  2983 => x"000034d2",
  2984 => x"0000201e",
  2985 => x"00000002",
  2986 => x"000034f0",
  2987 => x"0000201e",
  2988 => x"00000004",
  2989 => x"000029c4",
  2990 => x"00000000",
  2991 => x"00000000",
  2992 => x"00000000",
  2993 => x"000021f9",
  2994 => x"00000000",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memAWriteEnable = '1') and (from_zpu.memBWriteEnable = '1') and (from_zpu.memAAddr=from_zpu.memBAddr) and (from_zpu.memAWrite/=from_zpu.memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (from_zpu.memAWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memAWrite;
			to_zpu.memARead <= from_zpu.memAWrite;
		else
			to_zpu.memARead <= ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memBWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memBWrite;
			to_zpu.memBRead <= from_zpu.memBWrite;
		else
			to_zpu.memBRead <= ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;


end arch;

