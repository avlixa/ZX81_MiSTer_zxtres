-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Alastair M. Robinson for the ZPUFlex project.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.zpupkg.all;

entity CtrlROM_ROM is
generic
	(
		maxAddrBitBRAM : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_zpu : in ZPU_ToROM;
	to_zpu : out ZPU_FromROM
);
end CtrlROM_ROM;

architecture arch of CtrlROM_ROM is

type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"0b0b0b0b",
     1 => x"8c0b0b0b",
     2 => x"0b81e004",
     3 => x"0b0b0b0b",
     4 => x"8c04ff0d",
     5 => x"80040400",
     6 => x"00000016",
     7 => x"00000000",
     8 => x"0b0b80d1",
     9 => x"c4080b0b",
    10 => x"80d1c808",
    11 => x"0b0b80d1",
    12 => x"cc080b0b",
    13 => x"0b0b9808",
    14 => x"2d0b0b80",
    15 => x"d1cc0c0b",
    16 => x"0b80d1c8",
    17 => x"0c0b0b80",
    18 => x"d1c40c04",
    19 => x"00000000",
    20 => x"00000000",
    21 => x"00000000",
    22 => x"00000000",
    23 => x"00000000",
    24 => x"71fd0608",
    25 => x"72830609",
    26 => x"81058205",
    27 => x"832b2a83",
    28 => x"ffff0652",
    29 => x"0471fc06",
    30 => x"08728306",
    31 => x"09810583",
    32 => x"05101010",
    33 => x"2a81ff06",
    34 => x"520471fd",
    35 => x"060883ff",
    36 => x"ff738306",
    37 => x"09810582",
    38 => x"05832b2b",
    39 => x"09067383",
    40 => x"ffff0673",
    41 => x"83060981",
    42 => x"05820583",
    43 => x"2b0b2b07",
    44 => x"72fc060c",
    45 => x"51510471",
    46 => x"fc06080b",
    47 => x"0b0bbdc0",
    48 => x"73830610",
    49 => x"10050806",
    50 => x"7381ff06",
    51 => x"73830609",
    52 => x"81058305",
    53 => x"1010102b",
    54 => x"0772fc06",
    55 => x"0c515104",
    56 => x"80d1c470",
    57 => x"80dc8027",
    58 => x"8b388071",
    59 => x"70840553",
    60 => x"0c81e304",
    61 => x"8c518aa2",
    62 => x"0402fc05",
    63 => x"0df88051",
    64 => x"8f0b80d1",
    65 => x"d40c9f0b",
    66 => x"80d1d80c",
    67 => x"a0717081",
    68 => x"05533480",
    69 => x"d1d808ff",
    70 => x"0580d1d8",
    71 => x"0c80d1d8",
    72 => x"088025e8",
    73 => x"3880d1d4",
    74 => x"08ff0580",
    75 => x"d1d40c80",
    76 => x"d1d40880",
    77 => x"25d03880",
    78 => x"0b80d1d8",
    79 => x"0c800b80",
    80 => x"d1d40c02",
    81 => x"84050d04",
    82 => x"02f0050d",
    83 => x"f88053f8",
    84 => x"a05483bf",
    85 => x"52737081",
    86 => x"05553351",
    87 => x"70737081",
    88 => x"055534ff",
    89 => x"12527180",
    90 => x"25eb38fb",
    91 => x"c0539f52",
    92 => x"a0737081",
    93 => x"055534ff",
    94 => x"12527180",
    95 => x"25f23802",
    96 => x"90050d04",
    97 => x"02f4050d",
    98 => x"74538e0b",
    99 => x"80d1d408",
   100 => x"25913882",
   101 => x"c82d80d1",
   102 => x"d408ff05",
   103 => x"80d1d40c",
   104 => x"838a0480",
   105 => x"d1d40880",
   106 => x"d1d80853",
   107 => x"51728a2e",
   108 => x"098106be",
   109 => x"38715171",
   110 => x"9f24a438",
   111 => x"80d1d408",
   112 => x"a02911f8",
   113 => x"80115151",
   114 => x"a0713480",
   115 => x"d1d80881",
   116 => x"0580d1d8",
   117 => x"0c80d1d8",
   118 => x"08519f71",
   119 => x"25de3880",
   120 => x"0b80d1d8",
   121 => x"0c80d1d4",
   122 => x"08810580",
   123 => x"d1d40c84",
   124 => x"880470a0",
   125 => x"2912f880",
   126 => x"11515172",
   127 => x"713480d1",
   128 => x"d8088105",
   129 => x"80d1d80c",
   130 => x"80d1d808",
   131 => x"a02e0981",
   132 => x"06913880",
   133 => x"0b80d1d8",
   134 => x"0c80d1d4",
   135 => x"08810580",
   136 => x"d1d40c02",
   137 => x"8c050d04",
   138 => x"02e8050d",
   139 => x"77795656",
   140 => x"880bfc16",
   141 => x"77712c8f",
   142 => x"06545254",
   143 => x"80537272",
   144 => x"25953871",
   145 => x"53fbe014",
   146 => x"51877134",
   147 => x"8114ff14",
   148 => x"545472f1",
   149 => x"387153f9",
   150 => x"1576712c",
   151 => x"87065351",
   152 => x"71802e8b",
   153 => x"38fbe014",
   154 => x"51717134",
   155 => x"81145472",
   156 => x"8e249538",
   157 => x"8f733153",
   158 => x"fbe01451",
   159 => x"a0713481",
   160 => x"14ff1454",
   161 => x"5472f138",
   162 => x"0298050d",
   163 => x"0402ec05",
   164 => x"0d800b80",
   165 => x"d1dc0cf6",
   166 => x"8c08f690",
   167 => x"0871882c",
   168 => x"565381ff",
   169 => x"06537373",
   170 => x"25893872",
   171 => x"54820b80",
   172 => x"d1dc0c71",
   173 => x"882c7281",
   174 => x"ff065355",
   175 => x"7472258d",
   176 => x"387180d1",
   177 => x"dc088407",
   178 => x"80d1dc0c",
   179 => x"5573842b",
   180 => x"75832b56",
   181 => x"5485bc74",
   182 => x"258f3882",
   183 => x"0b0b0b80",
   184 => x"c8fc0c80",
   185 => x"d05385f3",
   186 => x"04810b0b",
   187 => x"0b80c8fc",
   188 => x"0cbc530b",
   189 => x"0b80c8fc",
   190 => x"0881712b",
   191 => x"ff05f688",
   192 => x"0cfc0875",
   193 => x"7531ffb0",
   194 => x"05ff1371",
   195 => x"712cff94",
   196 => x"1a709f2a",
   197 => x"1170812c",
   198 => x"80d1dc08",
   199 => x"52545153",
   200 => x"57535152",
   201 => x"5276802e",
   202 => x"85387081",
   203 => x"075170f6",
   204 => x"940c7209",
   205 => x"8105f680",
   206 => x"0c710981",
   207 => x"05f6840c",
   208 => x"0294050d",
   209 => x"0402f405",
   210 => x"0d745372",
   211 => x"70810554",
   212 => x"80f52d52",
   213 => x"71802e89",
   214 => x"38715183",
   215 => x"842d86cb",
   216 => x"04810b80",
   217 => x"d1c40c02",
   218 => x"8c050d04",
   219 => x"02fc050d",
   220 => x"81808051",
   221 => x"c0115170",
   222 => x"fb380284",
   223 => x"050d0402",
   224 => x"fc050dec",
   225 => x"5183710c",
   226 => x"86ec2d82",
   227 => x"710c0284",
   228 => x"050d0402",
   229 => x"fc050d84",
   230 => x"bf5186ec",
   231 => x"2dff1151",
   232 => x"708025f6",
   233 => x"38028405",
   234 => x"0d040402",
   235 => x"fc050d92",
   236 => x"ce2d80d1",
   237 => x"c40880cf",
   238 => x"800c80cd",
   239 => x"dc519586",
   240 => x"2d028405",
   241 => x"0d0402fc",
   242 => x"050d92ce",
   243 => x"2d80d1c4",
   244 => x"0880cdcc",
   245 => x"0c80cca8",
   246 => x"5195862d",
   247 => x"0284050d",
   248 => x"0402dc05",
   249 => x"0d7a5580",
   250 => x"59840bec",
   251 => x"0c80c984",
   252 => x"085380c9",
   253 => x"8008812e",
   254 => x"0981068c",
   255 => x"38728280",
   256 => x"0780c984",
   257 => x"0c889304",
   258 => x"72828007",
   259 => x"82803280",
   260 => x"c9840c80",
   261 => x"c98408fc",
   262 => x"0c86ec2d",
   263 => x"745280d1",
   264 => x"e051b3fd",
   265 => x"2d80d1c4",
   266 => x"08802e81",
   267 => x"ae3880d1",
   268 => x"e4085480",
   269 => x"5673852e",
   270 => x"098106a5",
   271 => x"38745186",
   272 => x"c52d8793",
   273 => x"2d87932d",
   274 => x"87932d87",
   275 => x"932d8793",
   276 => x"2d87932d",
   277 => x"80d1ec08",
   278 => x"5195862d",
   279 => x"81538a98",
   280 => x"0473f80c",
   281 => x"a50bec0c",
   282 => x"87932d84",
   283 => x"0bec0c75",
   284 => x"ff155758",
   285 => x"75802e8b",
   286 => x"38811876",
   287 => x"812a5758",
   288 => x"88f404f7",
   289 => x"18588159",
   290 => x"80742580",
   291 => x"ce387752",
   292 => x"755184a8",
   293 => x"2d80d2b8",
   294 => x"5280d1e0",
   295 => x"51b6ca2d",
   296 => x"80d1c408",
   297 => x"802e9b38",
   298 => x"80d2b857",
   299 => x"83fc5576",
   300 => x"70840558",
   301 => x"08e80cfc",
   302 => x"15557480",
   303 => x"25f13889",
   304 => x"ca0480d1",
   305 => x"c4085984",
   306 => x"805480d1",
   307 => x"e051b69a",
   308 => x"2dfc8014",
   309 => x"81175754",
   310 => x"89880480",
   311 => x"c9800853",
   312 => x"72893872",
   313 => x"5186ff2d",
   314 => x"8a820480",
   315 => x"0b80c980",
   316 => x"0c80c984",
   317 => x"08828007",
   318 => x"82803270",
   319 => x"80c9840c",
   320 => x"fc0c7880",
   321 => x"2e893880",
   322 => x"d1ec0851",
   323 => x"8a930480",
   324 => x"cc845195",
   325 => x"862d7853",
   326 => x"7280d1c4",
   327 => x"0c02a405",
   328 => x"0d0402e4",
   329 => x"050d900b",
   330 => x"80c9840c",
   331 => x"805186ff",
   332 => x"2d805186",
   333 => x"ff2d840b",
   334 => x"ec0c929e",
   335 => x"2d8ec92d",
   336 => x"81f92d83",
   337 => x"5392812d",
   338 => x"8151858d",
   339 => x"2dff1353",
   340 => x"728025f1",
   341 => x"38840bec",
   342 => x"0c80c7b0",
   343 => x"5186c52d",
   344 => x"aab52d80",
   345 => x"d1c40880",
   346 => x"2e83c738",
   347 => x"810bec0c",
   348 => x"840bec0c",
   349 => x"bdd05280",
   350 => x"d1e051b3",
   351 => x"fd2d80d1",
   352 => x"c408802e",
   353 => x"80cb3880",
   354 => x"d2b85280",
   355 => x"d1e051b6",
   356 => x"ca2d80d1",
   357 => x"c408802e",
   358 => x"b83880d2",
   359 => x"b80b80f5",
   360 => x"2d80cff0",
   361 => x"0c80d2b9",
   362 => x"0b80f52d",
   363 => x"80cff40c",
   364 => x"80d2ba0b",
   365 => x"80f52d80",
   366 => x"cff80c80",
   367 => x"d2bb0b80",
   368 => x"f52d80cf",
   369 => x"fc0c80d2",
   370 => x"bc0b80f5",
   371 => x"2d80d080",
   372 => x"0cbde052",
   373 => x"80d1e051",
   374 => x"b3fd2d80",
   375 => x"d1c40880",
   376 => x"2e80cb38",
   377 => x"80d2b852",
   378 => x"80d1e051",
   379 => x"b6ca2d80",
   380 => x"d1c40880",
   381 => x"2eb83880",
   382 => x"d2b80b80",
   383 => x"f52d80cf",
   384 => x"dc0c80d2",
   385 => x"b90b80f5",
   386 => x"2d80cfe0",
   387 => x"0c80d2ba",
   388 => x"0b80f52d",
   389 => x"80cfe40c",
   390 => x"80d2bb0b",
   391 => x"80f52d80",
   392 => x"cfe80c80",
   393 => x"d2bc0b80",
   394 => x"f52d80cf",
   395 => x"ec0c87e1",
   396 => x"51bdba2d",
   397 => x"80c98408",
   398 => x"80cfd80c",
   399 => x"80c98408",
   400 => x"fc0c80d2",
   401 => x"9808882a",
   402 => x"70810651",
   403 => x"5372802e",
   404 => x"8c3880ca",
   405 => x"d00b80d1",
   406 => x"ec0c8ce5",
   407 => x"0480c988",
   408 => x"0b80d1ec",
   409 => x"0c80d1ec",
   410 => x"08519586",
   411 => x"2d860b80",
   412 => x"d2ac0c92",
   413 => x"d72d8ed5",
   414 => x"2d95992d",
   415 => x"80d1c408",
   416 => x"80d1ec08",
   417 => x"80e81180",
   418 => x"f52d7084",
   419 => x"2b7080c9",
   420 => x"840c80f4",
   421 => x"1380f52d",
   422 => x"70852b72",
   423 => x"077080c9",
   424 => x"840c80d2",
   425 => x"9808882a",
   426 => x"70810681",
   427 => x"801780f5",
   428 => x"2d80cfd8",
   429 => x"08555751",
   430 => x"53535a56",
   431 => x"57555772",
   432 => x"802e8b38",
   433 => x"73822b87",
   434 => x"fc06538d",
   435 => x"d6047389",
   436 => x"2b87fc80",
   437 => x"06537473",
   438 => x"0780c984",
   439 => x"0c758106",
   440 => x"5372802e",
   441 => x"8b3880c9",
   442 => x"84088107",
   443 => x"80c9840c",
   444 => x"75812a70",
   445 => x"81065153",
   446 => x"72802e8b",
   447 => x"3880c984",
   448 => x"08820780",
   449 => x"c9840c75",
   450 => x"822a7081",
   451 => x"06515372",
   452 => x"802e8c38",
   453 => x"80c98408",
   454 => x"81800780",
   455 => x"c9840c80",
   456 => x"c98408fc",
   457 => x"0c865376",
   458 => x"83388453",
   459 => x"72ec0c8c",
   460 => x"f604800b",
   461 => x"80d1c40c",
   462 => x"029c050d",
   463 => x"0471980c",
   464 => x"04ffb008",
   465 => x"80d1c40c",
   466 => x"04810bff",
   467 => x"b00c0480",
   468 => x"0bffb00c",
   469 => x"0402f405",
   470 => x"0d8fe304",
   471 => x"80d1c408",
   472 => x"81f02e09",
   473 => x"81068a38",
   474 => x"810b80cf",
   475 => x"d00c8fe3",
   476 => x"0480d1c4",
   477 => x"0881e02e",
   478 => x"0981068a",
   479 => x"38810b80",
   480 => x"cfd40c8f",
   481 => x"e30480d1",
   482 => x"c4085280",
   483 => x"cfd40880",
   484 => x"2e893880",
   485 => x"d1c40881",
   486 => x"80055271",
   487 => x"842c728f",
   488 => x"06535380",
   489 => x"cfd00880",
   490 => x"2e9a3872",
   491 => x"842980cf",
   492 => x"90057213",
   493 => x"81712b70",
   494 => x"09730806",
   495 => x"730c5153",
   496 => x"538fd704",
   497 => x"72842980",
   498 => x"cf900572",
   499 => x"1383712b",
   500 => x"72080772",
   501 => x"0c535380",
   502 => x"0b80cfd4",
   503 => x"0c800b80",
   504 => x"cfd00c80",
   505 => x"d1f05190",
   506 => x"ea2d80d1",
   507 => x"c408ff24",
   508 => x"feea3880",
   509 => x"0b80d1c4",
   510 => x"0c028c05",
   511 => x"0d0402f8",
   512 => x"050d80cf",
   513 => x"90528f51",
   514 => x"80727084",
   515 => x"05540cff",
   516 => x"11517080",
   517 => x"25f23802",
   518 => x"88050d04",
   519 => x"02f0050d",
   520 => x"75518ecf",
   521 => x"2d70822c",
   522 => x"fc0680cf",
   523 => x"90117210",
   524 => x"9e067108",
   525 => x"70722a70",
   526 => x"83068274",
   527 => x"2b700974",
   528 => x"06760c54",
   529 => x"51565753",
   530 => x"51538ec9",
   531 => x"2d7180d1",
   532 => x"c40c0290",
   533 => x"050d0402",
   534 => x"fc050d72",
   535 => x"5180710c",
   536 => x"800b8412",
   537 => x"0c028405",
   538 => x"0d0402f0",
   539 => x"050d7570",
   540 => x"08841208",
   541 => x"535353ff",
   542 => x"5471712e",
   543 => x"a8388ecf",
   544 => x"2d841308",
   545 => x"70842914",
   546 => x"88117008",
   547 => x"7081ff06",
   548 => x"84180881",
   549 => x"11870684",
   550 => x"1a0c5351",
   551 => x"55515151",
   552 => x"8ec92d71",
   553 => x"547380d1",
   554 => x"c40c0290",
   555 => x"050d0402",
   556 => x"f4050d8e",
   557 => x"cf2de008",
   558 => x"708b2a70",
   559 => x"81065152",
   560 => x"5370802e",
   561 => x"a13880d1",
   562 => x"f0087084",
   563 => x"2980d1f8",
   564 => x"057481ff",
   565 => x"06710c51",
   566 => x"5180d1f0",
   567 => x"08811187",
   568 => x"0680d1f0",
   569 => x"0c51728c",
   570 => x"2c83ff06",
   571 => x"80d2980c",
   572 => x"800b80d2",
   573 => x"9c0c8ec1",
   574 => x"2d8ec92d",
   575 => x"028c050d",
   576 => x"0402fc05",
   577 => x"0d8ecf2d",
   578 => x"810b80d2",
   579 => x"9c0c8ec9",
   580 => x"2d80d29c",
   581 => x"085170f9",
   582 => x"38028405",
   583 => x"0d0402fc",
   584 => x"050d80d1",
   585 => x"f05190d7",
   586 => x"2d8ffe2d",
   587 => x"91af518e",
   588 => x"bd2d0284",
   589 => x"050d0402",
   590 => x"fc050d8f",
   591 => x"cf5186ec",
   592 => x"2dff1151",
   593 => x"708025f6",
   594 => x"38028405",
   595 => x"0d0480d2",
   596 => x"a40880d1",
   597 => x"c40c0402",
   598 => x"fc050d81",
   599 => x"0b80d084",
   600 => x"0c815185",
   601 => x"8d2d0284",
   602 => x"050d0402",
   603 => x"fc050d92",
   604 => x"f5048ed5",
   605 => x"2d80f651",
   606 => x"909c2d80",
   607 => x"d1c408f2",
   608 => x"3880da51",
   609 => x"909c2d80",
   610 => x"d1c408e6",
   611 => x"3880d080",
   612 => x"0851909c",
   613 => x"2d80d1c4",
   614 => x"08d83880",
   615 => x"d1c40880",
   616 => x"d0840c80",
   617 => x"d1c40851",
   618 => x"858d2d02",
   619 => x"84050d04",
   620 => x"02ec050d",
   621 => x"76548052",
   622 => x"870b8815",
   623 => x"80f52d56",
   624 => x"53747224",
   625 => x"8338a053",
   626 => x"72518384",
   627 => x"2d81128b",
   628 => x"1580f52d",
   629 => x"54527272",
   630 => x"25de3802",
   631 => x"94050d04",
   632 => x"02f0050d",
   633 => x"80d2a408",
   634 => x"5481f92d",
   635 => x"800b80d2",
   636 => x"a80c7308",
   637 => x"802e8189",
   638 => x"38820b80",
   639 => x"d1d80c80",
   640 => x"d2a8088f",
   641 => x"0680d1d4",
   642 => x"0c730852",
   643 => x"71832e96",
   644 => x"38718326",
   645 => x"89387181",
   646 => x"2eb03894",
   647 => x"ea047185",
   648 => x"2ea03894",
   649 => x"ea048814",
   650 => x"80f52d84",
   651 => x"150880c7",
   652 => x"c8535452",
   653 => x"86c52d71",
   654 => x"84291370",
   655 => x"08525294",
   656 => x"ee047351",
   657 => x"93b02d94",
   658 => x"ea0480cf",
   659 => x"d8088815",
   660 => x"082c7081",
   661 => x"06515271",
   662 => x"802e8838",
   663 => x"80c7cc51",
   664 => x"94e70480",
   665 => x"c7d05186",
   666 => x"c52d8414",
   667 => x"085186c5",
   668 => x"2d80d2a8",
   669 => x"08810580",
   670 => x"d2a80c8c",
   671 => x"145493f2",
   672 => x"04029005",
   673 => x"0d047180",
   674 => x"d2a40c93",
   675 => x"e02d80d2",
   676 => x"a808ff05",
   677 => x"80d2ac0c",
   678 => x"0402e805",
   679 => x"0d80d2a4",
   680 => x"0880d2b0",
   681 => x"08575580",
   682 => x"f651909c",
   683 => x"2d80d1c4",
   684 => x"08812a70",
   685 => x"81065152",
   686 => x"71802ea2",
   687 => x"3895c304",
   688 => x"8ed52d80",
   689 => x"f651909c",
   690 => x"2d80d1c4",
   691 => x"08f23880",
   692 => x"d0840881",
   693 => x"327080d0",
   694 => x"840c5185",
   695 => x"8d2d800b",
   696 => x"80d2a00c",
   697 => x"8651909c",
   698 => x"2d80d1c4",
   699 => x"08812a70",
   700 => x"81065152",
   701 => x"71802e8b",
   702 => x"3880c984",
   703 => x"08903280",
   704 => x"c9840c8c",
   705 => x"51909c2d",
   706 => x"80d1c408",
   707 => x"812a7081",
   708 => x"06515271",
   709 => x"802e80d1",
   710 => x"3880cfdc",
   711 => x"0880cff0",
   712 => x"0880cfdc",
   713 => x"0c80cff0",
   714 => x"0c80cfe0",
   715 => x"0880cff4",
   716 => x"0880cfe0",
   717 => x"0c80cff4",
   718 => x"0c80cfe4",
   719 => x"0880cff8",
   720 => x"0880cfe4",
   721 => x"0c80cff8",
   722 => x"0c80cfe8",
   723 => x"0880cffc",
   724 => x"0880cfe8",
   725 => x"0c80cffc",
   726 => x"0c80cfec",
   727 => x"0880d080",
   728 => x"0880cfec",
   729 => x"0c80d080",
   730 => x"0c80d298",
   731 => x"08a00652",
   732 => x"80722596",
   733 => x"3892b72d",
   734 => x"8ed52d80",
   735 => x"d0840881",
   736 => x"327080d0",
   737 => x"840c5185",
   738 => x"8d2d80d0",
   739 => x"840882ef",
   740 => x"3880cff0",
   741 => x"0851909c",
   742 => x"2d80d1c4",
   743 => x"08802e8b",
   744 => x"3880d2a0",
   745 => x"08810780",
   746 => x"d2a00c80",
   747 => x"cff40851",
   748 => x"909c2d80",
   749 => x"d1c40880",
   750 => x"2e8b3880",
   751 => x"d2a00882",
   752 => x"0780d2a0",
   753 => x"0c80cff8",
   754 => x"0851909c",
   755 => x"2d80d1c4",
   756 => x"08802e8b",
   757 => x"3880d2a0",
   758 => x"08840780",
   759 => x"d2a00c80",
   760 => x"cffc0851",
   761 => x"909c2d80",
   762 => x"d1c40880",
   763 => x"2e8b3880",
   764 => x"d2a00888",
   765 => x"0780d2a0",
   766 => x"0c80d080",
   767 => x"0851909c",
   768 => x"2d80d1c4",
   769 => x"08802e8b",
   770 => x"3880d2a0",
   771 => x"08900780",
   772 => x"d2a00c80",
   773 => x"cfdc0851",
   774 => x"909c2d80",
   775 => x"d1c40880",
   776 => x"2e8c3880",
   777 => x"d2a00882",
   778 => x"800780d2",
   779 => x"a00c80cf",
   780 => x"e0085190",
   781 => x"9c2d80d1",
   782 => x"c408802e",
   783 => x"8c3880d2",
   784 => x"a0088480",
   785 => x"0780d2a0",
   786 => x"0c80cfe4",
   787 => x"0851909c",
   788 => x"2d80d1c4",
   789 => x"08802e8c",
   790 => x"3880d2a0",
   791 => x"08888007",
   792 => x"80d2a00c",
   793 => x"80cfe808",
   794 => x"51909c2d",
   795 => x"80d1c408",
   796 => x"802e8c38",
   797 => x"80d2a008",
   798 => x"90800780",
   799 => x"d2a00c80",
   800 => x"cfec0851",
   801 => x"909c2d80",
   802 => x"d1c40880",
   803 => x"2e8c3880",
   804 => x"d2a008a0",
   805 => x"800780d2",
   806 => x"a00c9451",
   807 => x"909c2d80",
   808 => x"d1c40852",
   809 => x"9151909c",
   810 => x"2d7180d1",
   811 => x"c4080652",
   812 => x"80e65190",
   813 => x"9c2d7180",
   814 => x"d1c40806",
   815 => x"5271802e",
   816 => x"8d3880d2",
   817 => x"a0088480",
   818 => x"800780d2",
   819 => x"a00c80fe",
   820 => x"51909c2d",
   821 => x"80d1c408",
   822 => x"52875190",
   823 => x"9c2d7180",
   824 => x"d1c40807",
   825 => x"5271802e",
   826 => x"8d3880d2",
   827 => x"a0088880",
   828 => x"800780d2",
   829 => x"a00c80d2",
   830 => x"a008ed0c",
   831 => x"a28a0494",
   832 => x"51909c2d",
   833 => x"80d1c408",
   834 => x"52915190",
   835 => x"9c2d7180",
   836 => x"d1c40806",
   837 => x"5280e651",
   838 => x"909c2d71",
   839 => x"80d1c408",
   840 => x"06527180",
   841 => x"2e8d3880",
   842 => x"d2a00884",
   843 => x"80800780",
   844 => x"d2a00c80",
   845 => x"fe51909c",
   846 => x"2d80d1c4",
   847 => x"08528751",
   848 => x"909c2d71",
   849 => x"80d1c408",
   850 => x"07527180",
   851 => x"2e8d3880",
   852 => x"d2a00888",
   853 => x"80800780",
   854 => x"d2a00c80",
   855 => x"d2a008ed",
   856 => x"0c81f551",
   857 => x"909c2d80",
   858 => x"d1c40881",
   859 => x"2a708106",
   860 => x"515271a4",
   861 => x"3880cff0",
   862 => x"0851909c",
   863 => x"2d80d1c4",
   864 => x"08812a70",
   865 => x"81065152",
   866 => x"718e3880",
   867 => x"d2980881",
   868 => x"06528072",
   869 => x"2580c238",
   870 => x"80d29808",
   871 => x"81065280",
   872 => x"72258438",
   873 => x"92b72d80",
   874 => x"d2ac0852",
   875 => x"71802e8a",
   876 => x"38ff1280",
   877 => x"d2ac0c9b",
   878 => x"d90480d2",
   879 => x"a8081080",
   880 => x"d2a80805",
   881 => x"70842916",
   882 => x"51528812",
   883 => x"08802e89",
   884 => x"38ff5188",
   885 => x"12085271",
   886 => x"2d81f251",
   887 => x"909c2d80",
   888 => x"d1c40881",
   889 => x"2a708106",
   890 => x"515271a4",
   891 => x"3880cff4",
   892 => x"0851909c",
   893 => x"2d80d1c4",
   894 => x"08812a70",
   895 => x"81065152",
   896 => x"718e3880",
   897 => x"d2980882",
   898 => x"06528072",
   899 => x"2580c338",
   900 => x"80d29808",
   901 => x"82065280",
   902 => x"72258438",
   903 => x"92b72d80",
   904 => x"d2a808ff",
   905 => x"1180d2ac",
   906 => x"08565353",
   907 => x"7372258a",
   908 => x"38811480",
   909 => x"d2ac0c9c",
   910 => x"d2047210",
   911 => x"13708429",
   912 => x"16515288",
   913 => x"1208802e",
   914 => x"8938fe51",
   915 => x"88120852",
   916 => x"712d81fd",
   917 => x"51909c2d",
   918 => x"80d1c408",
   919 => x"812a7081",
   920 => x"06515271",
   921 => x"a43880cf",
   922 => x"f8085190",
   923 => x"9c2d80d1",
   924 => x"c408812a",
   925 => x"70810651",
   926 => x"52718e38",
   927 => x"80d29808",
   928 => x"84065280",
   929 => x"722580c0",
   930 => x"3880d298",
   931 => x"08840652",
   932 => x"80722584",
   933 => x"3892b72d",
   934 => x"80d2ac08",
   935 => x"802e8a38",
   936 => x"800b80d2",
   937 => x"ac0c9dc8",
   938 => x"0480d2a8",
   939 => x"081080d2",
   940 => x"a8080570",
   941 => x"84291651",
   942 => x"52881208",
   943 => x"802e8938",
   944 => x"fd518812",
   945 => x"0852712d",
   946 => x"81fa5190",
   947 => x"9c2d80d1",
   948 => x"c408812a",
   949 => x"70810651",
   950 => x"5271a438",
   951 => x"80cffc08",
   952 => x"51909c2d",
   953 => x"80d1c408",
   954 => x"812a7081",
   955 => x"06515271",
   956 => x"8e3880d2",
   957 => x"98088806",
   958 => x"52807225",
   959 => x"80c03880",
   960 => x"d2980888",
   961 => x"06528072",
   962 => x"25843892",
   963 => x"b72d80d2",
   964 => x"a808ff11",
   965 => x"545280d2",
   966 => x"ac087325",
   967 => x"89387280",
   968 => x"d2ac0c9e",
   969 => x"be047110",
   970 => x"12708429",
   971 => x"16515288",
   972 => x"1208802e",
   973 => x"8938fc51",
   974 => x"88120852",
   975 => x"712d80d2",
   976 => x"ac087053",
   977 => x"5473802e",
   978 => x"8a388c15",
   979 => x"ff155555",
   980 => x"9ec50482",
   981 => x"0b80d1d8",
   982 => x"0c718f06",
   983 => x"80d1d40c",
   984 => x"81eb5190",
   985 => x"9c2d80d1",
   986 => x"c408812a",
   987 => x"70810651",
   988 => x"5271802e",
   989 => x"ad387408",
   990 => x"852e0981",
   991 => x"06a43888",
   992 => x"1580f52d",
   993 => x"ff055271",
   994 => x"881681b7",
   995 => x"2d71982b",
   996 => x"52718025",
   997 => x"8838800b",
   998 => x"881681b7",
   999 => x"2d745193",
  1000 => x"b02d81f4",
  1001 => x"51909c2d",
  1002 => x"80d1c408",
  1003 => x"812a7081",
  1004 => x"06515271",
  1005 => x"802eb338",
  1006 => x"7408852e",
  1007 => x"098106aa",
  1008 => x"38881580",
  1009 => x"f52d8105",
  1010 => x"52718816",
  1011 => x"81b72d71",
  1012 => x"81ff068b",
  1013 => x"1680f52d",
  1014 => x"54527272",
  1015 => x"27873872",
  1016 => x"881681b7",
  1017 => x"2d745193",
  1018 => x"b02d80da",
  1019 => x"51909c2d",
  1020 => x"80d1c408",
  1021 => x"812a7081",
  1022 => x"06515271",
  1023 => x"8e3880d2",
  1024 => x"98089006",
  1025 => x"52807225",
  1026 => x"81bc3880",
  1027 => x"d2a40880",
  1028 => x"d2980890",
  1029 => x"06535380",
  1030 => x"72258438",
  1031 => x"92b72d80",
  1032 => x"d2ac0854",
  1033 => x"73802e8a",
  1034 => x"388c13ff",
  1035 => x"155553a0",
  1036 => x"a4047208",
  1037 => x"5271822e",
  1038 => x"a6387182",
  1039 => x"26893871",
  1040 => x"812eaa38",
  1041 => x"a1c60471",
  1042 => x"832eb438",
  1043 => x"71842e09",
  1044 => x"810680f2",
  1045 => x"38881308",
  1046 => x"5195862d",
  1047 => x"a1c60480",
  1048 => x"d2ac0851",
  1049 => x"88130852",
  1050 => x"712da1c6",
  1051 => x"04810b88",
  1052 => x"14082b80",
  1053 => x"cfd80832",
  1054 => x"80cfd80c",
  1055 => x"a19a0488",
  1056 => x"1380f52d",
  1057 => x"81058b14",
  1058 => x"80f52d53",
  1059 => x"54717424",
  1060 => x"83388054",
  1061 => x"73881481",
  1062 => x"b72d93e0",
  1063 => x"2da1c604",
  1064 => x"7508802e",
  1065 => x"a4387508",
  1066 => x"51909c2d",
  1067 => x"80d1c408",
  1068 => x"81065271",
  1069 => x"802e8c38",
  1070 => x"80d2ac08",
  1071 => x"51841608",
  1072 => x"52712d88",
  1073 => x"165675d8",
  1074 => x"38805480",
  1075 => x"0b80d1d8",
  1076 => x"0c738f06",
  1077 => x"80d1d40c",
  1078 => x"a0527380",
  1079 => x"d2ac082e",
  1080 => x"09810699",
  1081 => x"3880d2a8",
  1082 => x"08ff0574",
  1083 => x"32700981",
  1084 => x"05707207",
  1085 => x"9f2a9171",
  1086 => x"31515153",
  1087 => x"53715183",
  1088 => x"842d8114",
  1089 => x"548e7425",
  1090 => x"c23880d0",
  1091 => x"840880d1",
  1092 => x"c40c0298",
  1093 => x"050d0402",
  1094 => x"f4050dd4",
  1095 => x"5281ff72",
  1096 => x"0c710853",
  1097 => x"81ff720c",
  1098 => x"72882b83",
  1099 => x"fe800672",
  1100 => x"087081ff",
  1101 => x"06515253",
  1102 => x"81ff720c",
  1103 => x"72710788",
  1104 => x"2b720870",
  1105 => x"81ff0651",
  1106 => x"525381ff",
  1107 => x"720c7271",
  1108 => x"07882b72",
  1109 => x"087081ff",
  1110 => x"06720780",
  1111 => x"d1c40c52",
  1112 => x"53028c05",
  1113 => x"0d0402f4",
  1114 => x"050d7476",
  1115 => x"7181ff06",
  1116 => x"d40c5353",
  1117 => x"80d2b408",
  1118 => x"85387189",
  1119 => x"2b527198",
  1120 => x"2ad40c71",
  1121 => x"902a7081",
  1122 => x"ff06d40c",
  1123 => x"5171882a",
  1124 => x"7081ff06",
  1125 => x"d40c5171",
  1126 => x"81ff06d4",
  1127 => x"0c72902a",
  1128 => x"7081ff06",
  1129 => x"d40c51d4",
  1130 => x"087081ff",
  1131 => x"06515182",
  1132 => x"b8bf5270",
  1133 => x"81ff2e09",
  1134 => x"81069438",
  1135 => x"81ff0bd4",
  1136 => x"0cd40870",
  1137 => x"81ff06ff",
  1138 => x"14545151",
  1139 => x"71e53870",
  1140 => x"80d1c40c",
  1141 => x"028c050d",
  1142 => x"0402fc05",
  1143 => x"0d81c751",
  1144 => x"81ff0bd4",
  1145 => x"0cff1151",
  1146 => x"708025f4",
  1147 => x"38028405",
  1148 => x"0d0402f4",
  1149 => x"050d81ff",
  1150 => x"0bd40c93",
  1151 => x"53805287",
  1152 => x"fc80c151",
  1153 => x"a2e62d80",
  1154 => x"d1c4088b",
  1155 => x"3881ff0b",
  1156 => x"d40c8153",
  1157 => x"a4a004a3",
  1158 => x"d92dff13",
  1159 => x"5372de38",
  1160 => x"7280d1c4",
  1161 => x"0c028c05",
  1162 => x"0d0402ec",
  1163 => x"050d810b",
  1164 => x"80d2b40c",
  1165 => x"8454d008",
  1166 => x"708f2a70",
  1167 => x"81065151",
  1168 => x"5372f338",
  1169 => x"72d00ca3",
  1170 => x"d92d80c7",
  1171 => x"d45186c5",
  1172 => x"2dd00870",
  1173 => x"8f2a7081",
  1174 => x"06515153",
  1175 => x"72f33881",
  1176 => x"0bd00cb1",
  1177 => x"53805284",
  1178 => x"d480c051",
  1179 => x"a2e62d80",
  1180 => x"d1c40881",
  1181 => x"2e933872",
  1182 => x"822ebf38",
  1183 => x"ff135372",
  1184 => x"e438ff14",
  1185 => x"5473ffae",
  1186 => x"38a3d92d",
  1187 => x"83aa5284",
  1188 => x"9c80c851",
  1189 => x"a2e62d80",
  1190 => x"d1c40881",
  1191 => x"2e098106",
  1192 => x"9338a297",
  1193 => x"2d80d1c4",
  1194 => x"0883ffff",
  1195 => x"06537283",
  1196 => x"aa2e9f38",
  1197 => x"a3f22da5",
  1198 => x"cd0480c7",
  1199 => x"e05186c5",
  1200 => x"2d8053a7",
  1201 => x"a20480c7",
  1202 => x"f85186c5",
  1203 => x"2d8054a6",
  1204 => x"f30481ff",
  1205 => x"0bd40cb1",
  1206 => x"54a3d92d",
  1207 => x"8fcf5380",
  1208 => x"5287fc80",
  1209 => x"f751a2e6",
  1210 => x"2d80d1c4",
  1211 => x"085580d1",
  1212 => x"c408812e",
  1213 => x"0981069c",
  1214 => x"3881ff0b",
  1215 => x"d40c820a",
  1216 => x"52849c80",
  1217 => x"e951a2e6",
  1218 => x"2d80d1c4",
  1219 => x"08802e8d",
  1220 => x"38a3d92d",
  1221 => x"ff135372",
  1222 => x"c638a6e6",
  1223 => x"0481ff0b",
  1224 => x"d40c80d1",
  1225 => x"c4085287",
  1226 => x"fc80fa51",
  1227 => x"a2e62d80",
  1228 => x"d1c408b2",
  1229 => x"3881ff0b",
  1230 => x"d40cd408",
  1231 => x"5381ff0b",
  1232 => x"d40c81ff",
  1233 => x"0bd40c81",
  1234 => x"ff0bd40c",
  1235 => x"81ff0bd4",
  1236 => x"0c72862a",
  1237 => x"70810676",
  1238 => x"56515372",
  1239 => x"963880d1",
  1240 => x"c40854a6",
  1241 => x"f3047382",
  1242 => x"2efedb38",
  1243 => x"ff145473",
  1244 => x"fee73873",
  1245 => x"80d2b40c",
  1246 => x"738b3881",
  1247 => x"5287fc80",
  1248 => x"d051a2e6",
  1249 => x"2d81ff0b",
  1250 => x"d40cd008",
  1251 => x"708f2a70",
  1252 => x"81065151",
  1253 => x"5372f338",
  1254 => x"72d00c81",
  1255 => x"ff0bd40c",
  1256 => x"81537280",
  1257 => x"d1c40c02",
  1258 => x"94050d04",
  1259 => x"02e8050d",
  1260 => x"78558056",
  1261 => x"81ff0bd4",
  1262 => x"0cd00870",
  1263 => x"8f2a7081",
  1264 => x"06515153",
  1265 => x"72f33882",
  1266 => x"810bd00c",
  1267 => x"81ff0bd4",
  1268 => x"0c775287",
  1269 => x"fc80d151",
  1270 => x"a2e62d80",
  1271 => x"dbc6df54",
  1272 => x"80d1c408",
  1273 => x"802e8b38",
  1274 => x"80c89851",
  1275 => x"86c52da8",
  1276 => x"c60481ff",
  1277 => x"0bd40cd4",
  1278 => x"087081ff",
  1279 => x"06515372",
  1280 => x"81fe2e09",
  1281 => x"81069e38",
  1282 => x"80ff53a2",
  1283 => x"972d80d1",
  1284 => x"c4087570",
  1285 => x"8405570c",
  1286 => x"ff135372",
  1287 => x"8025ec38",
  1288 => x"8156a8ab",
  1289 => x"04ff1454",
  1290 => x"73c83881",
  1291 => x"ff0bd40c",
  1292 => x"81ff0bd4",
  1293 => x"0cd00870",
  1294 => x"8f2a7081",
  1295 => x"06515153",
  1296 => x"72f33872",
  1297 => x"d00c7580",
  1298 => x"d1c40c02",
  1299 => x"98050d04",
  1300 => x"02e8050d",
  1301 => x"77797b58",
  1302 => x"55558053",
  1303 => x"727625a3",
  1304 => x"38747081",
  1305 => x"055680f5",
  1306 => x"2d747081",
  1307 => x"055680f5",
  1308 => x"2d525271",
  1309 => x"712e8638",
  1310 => x"8151a985",
  1311 => x"04811353",
  1312 => x"a8dc0480",
  1313 => x"517080d1",
  1314 => x"c40c0298",
  1315 => x"050d0402",
  1316 => x"ec050d76",
  1317 => x"5574802e",
  1318 => x"80c2389a",
  1319 => x"1580e02d",
  1320 => x"51b7a42d",
  1321 => x"80d1c408",
  1322 => x"80d1c408",
  1323 => x"80d8e80c",
  1324 => x"80d1c408",
  1325 => x"545480d8",
  1326 => x"c408802e",
  1327 => x"9a389415",
  1328 => x"80e02d51",
  1329 => x"b7a42d80",
  1330 => x"d1c40890",
  1331 => x"2b83fff0",
  1332 => x"0a067075",
  1333 => x"07515372",
  1334 => x"80d8e80c",
  1335 => x"80d8e808",
  1336 => x"5372802e",
  1337 => x"9d3880d8",
  1338 => x"bc08fe14",
  1339 => x"712980d8",
  1340 => x"d0080580",
  1341 => x"d8ec0c70",
  1342 => x"842b80d8",
  1343 => x"c80c54aa",
  1344 => x"b00480d8",
  1345 => x"d40880d8",
  1346 => x"e80c80d8",
  1347 => x"d80880d8",
  1348 => x"ec0c80d8",
  1349 => x"c408802e",
  1350 => x"8b3880d8",
  1351 => x"bc08842b",
  1352 => x"53aaab04",
  1353 => x"80d8dc08",
  1354 => x"842b5372",
  1355 => x"80d8c80c",
  1356 => x"0294050d",
  1357 => x"0402d805",
  1358 => x"0d800b80",
  1359 => x"d8c40c84",
  1360 => x"54a4aa2d",
  1361 => x"80d1c408",
  1362 => x"802e9738",
  1363 => x"80d2b852",
  1364 => x"8051a7ac",
  1365 => x"2d80d1c4",
  1366 => x"08802e86",
  1367 => x"38fe54aa",
  1368 => x"ea04ff14",
  1369 => x"54738024",
  1370 => x"d838738d",
  1371 => x"3880c8a8",
  1372 => x"5186c52d",
  1373 => x"7355b0bf",
  1374 => x"04805681",
  1375 => x"0b80d8f0",
  1376 => x"0c885380",
  1377 => x"c8bc5280",
  1378 => x"d2ee51a8",
  1379 => x"d02d80d1",
  1380 => x"c408762e",
  1381 => x"09810689",
  1382 => x"3880d1c4",
  1383 => x"0880d8f0",
  1384 => x"0c885380",
  1385 => x"c8c85280",
  1386 => x"d38a51a8",
  1387 => x"d02d80d1",
  1388 => x"c4088938",
  1389 => x"80d1c408",
  1390 => x"80d8f00c",
  1391 => x"80d8f008",
  1392 => x"802e8181",
  1393 => x"3880d5fe",
  1394 => x"0b80f52d",
  1395 => x"80d5ff0b",
  1396 => x"80f52d71",
  1397 => x"982b7190",
  1398 => x"2b0780d6",
  1399 => x"800b80f5",
  1400 => x"2d70882b",
  1401 => x"720780d6",
  1402 => x"810b80f5",
  1403 => x"2d710780",
  1404 => x"d6b60b80",
  1405 => x"f52d80d6",
  1406 => x"b70b80f5",
  1407 => x"2d71882b",
  1408 => x"07535f54",
  1409 => x"525a5657",
  1410 => x"557381ab",
  1411 => x"aa2e0981",
  1412 => x"068e3875",
  1413 => x"51b6f32d",
  1414 => x"80d1c408",
  1415 => x"56acae04",
  1416 => x"7382d4d5",
  1417 => x"2e883880",
  1418 => x"c8d451ac",
  1419 => x"fa0480d2",
  1420 => x"b8527551",
  1421 => x"a7ac2d80",
  1422 => x"d1c40855",
  1423 => x"80d1c408",
  1424 => x"802e83fb",
  1425 => x"38885380",
  1426 => x"c8c85280",
  1427 => x"d38a51a8",
  1428 => x"d02d80d1",
  1429 => x"c4088a38",
  1430 => x"810b80d8",
  1431 => x"c40cad80",
  1432 => x"04885380",
  1433 => x"c8bc5280",
  1434 => x"d2ee51a8",
  1435 => x"d02d80d1",
  1436 => x"c408802e",
  1437 => x"8b3880c8",
  1438 => x"e85186c5",
  1439 => x"2daddf04",
  1440 => x"80d6b60b",
  1441 => x"80f52d54",
  1442 => x"7380d52e",
  1443 => x"09810680",
  1444 => x"ce3880d6",
  1445 => x"b70b80f5",
  1446 => x"2d547381",
  1447 => x"aa2e0981",
  1448 => x"06bd3880",
  1449 => x"0b80d2b8",
  1450 => x"0b80f52d",
  1451 => x"56547481",
  1452 => x"e92e8338",
  1453 => x"81547481",
  1454 => x"eb2e8c38",
  1455 => x"80557375",
  1456 => x"2e098106",
  1457 => x"82f93880",
  1458 => x"d2c30b80",
  1459 => x"f52d5574",
  1460 => x"8e3880d2",
  1461 => x"c40b80f5",
  1462 => x"2d547382",
  1463 => x"2e863880",
  1464 => x"55b0bf04",
  1465 => x"80d2c50b",
  1466 => x"80f52d70",
  1467 => x"80d8bc0c",
  1468 => x"ff0580d8",
  1469 => x"c00c80d2",
  1470 => x"c60b80f5",
  1471 => x"2d80d2c7",
  1472 => x"0b80f52d",
  1473 => x"58760577",
  1474 => x"82802905",
  1475 => x"7080d8cc",
  1476 => x"0c80d2c8",
  1477 => x"0b80f52d",
  1478 => x"7080d8e0",
  1479 => x"0c80d8c4",
  1480 => x"08595758",
  1481 => x"76802e81",
  1482 => x"b7388853",
  1483 => x"80c8c852",
  1484 => x"80d38a51",
  1485 => x"a8d02d80",
  1486 => x"d1c40882",
  1487 => x"823880d8",
  1488 => x"bc087084",
  1489 => x"2b80d8c8",
  1490 => x"0c7080d8",
  1491 => x"dc0c80d2",
  1492 => x"dd0b80f5",
  1493 => x"2d80d2dc",
  1494 => x"0b80f52d",
  1495 => x"71828029",
  1496 => x"0580d2de",
  1497 => x"0b80f52d",
  1498 => x"70848080",
  1499 => x"291280d2",
  1500 => x"df0b80f5",
  1501 => x"2d708180",
  1502 => x"0a291270",
  1503 => x"80d8e40c",
  1504 => x"80d8e008",
  1505 => x"712980d8",
  1506 => x"cc080570",
  1507 => x"80d8d00c",
  1508 => x"80d2e50b",
  1509 => x"80f52d80",
  1510 => x"d2e40b80",
  1511 => x"f52d7182",
  1512 => x"80290580",
  1513 => x"d2e60b80",
  1514 => x"f52d7084",
  1515 => x"80802912",
  1516 => x"80d2e70b",
  1517 => x"80f52d70",
  1518 => x"982b81f0",
  1519 => x"0a067205",
  1520 => x"7080d8d4",
  1521 => x"0cfe117e",
  1522 => x"29770580",
  1523 => x"d8d80c52",
  1524 => x"59524354",
  1525 => x"5e515259",
  1526 => x"525d5759",
  1527 => x"57b0b804",
  1528 => x"80d2ca0b",
  1529 => x"80f52d80",
  1530 => x"d2c90b80",
  1531 => x"f52d7182",
  1532 => x"80290570",
  1533 => x"80d8c80c",
  1534 => x"70a02983",
  1535 => x"ff057089",
  1536 => x"2a7080d8",
  1537 => x"dc0c80d2",
  1538 => x"cf0b80f5",
  1539 => x"2d80d2ce",
  1540 => x"0b80f52d",
  1541 => x"71828029",
  1542 => x"057080d8",
  1543 => x"e40c7b71",
  1544 => x"291e7080",
  1545 => x"d8d80c7d",
  1546 => x"80d8d40c",
  1547 => x"730580d8",
  1548 => x"d00c555e",
  1549 => x"51515555",
  1550 => x"8051a98f",
  1551 => x"2d815574",
  1552 => x"80d1c40c",
  1553 => x"02a8050d",
  1554 => x"0402ec05",
  1555 => x"0d767087",
  1556 => x"2c7180ff",
  1557 => x"06555654",
  1558 => x"80d8c408",
  1559 => x"8a387388",
  1560 => x"2c7481ff",
  1561 => x"06545580",
  1562 => x"d2b85280",
  1563 => x"d8cc0815",
  1564 => x"51a7ac2d",
  1565 => x"80d1c408",
  1566 => x"5480d1c4",
  1567 => x"08802eb8",
  1568 => x"3880d8c4",
  1569 => x"08802e9a",
  1570 => x"38728429",
  1571 => x"80d2b805",
  1572 => x"70085253",
  1573 => x"b6f32d80",
  1574 => x"d1c408f0",
  1575 => x"0a0653b1",
  1576 => x"b6047210",
  1577 => x"80d2b805",
  1578 => x"7080e02d",
  1579 => x"5253b7a4",
  1580 => x"2d80d1c4",
  1581 => x"08537254",
  1582 => x"7380d1c4",
  1583 => x"0c029405",
  1584 => x"0d0402e0",
  1585 => x"050d7970",
  1586 => x"842c80d8",
  1587 => x"ec080571",
  1588 => x"8f065255",
  1589 => x"53728a38",
  1590 => x"80d2b852",
  1591 => x"7351a7ac",
  1592 => x"2d72a029",
  1593 => x"80d2b805",
  1594 => x"54807480",
  1595 => x"f52d5653",
  1596 => x"74732e83",
  1597 => x"38815374",
  1598 => x"81e52e81",
  1599 => x"f4388170",
  1600 => x"74065458",
  1601 => x"72802e81",
  1602 => x"e8388b14",
  1603 => x"80f52d70",
  1604 => x"832a7906",
  1605 => x"5856769b",
  1606 => x"3880d088",
  1607 => x"08537289",
  1608 => x"387280d6",
  1609 => x"b80b81b7",
  1610 => x"2d7680d0",
  1611 => x"880c7353",
  1612 => x"b3f30475",
  1613 => x"8f2e0981",
  1614 => x"0681b638",
  1615 => x"749f068d",
  1616 => x"2980d6ab",
  1617 => x"11515381",
  1618 => x"1480f52d",
  1619 => x"73708105",
  1620 => x"5581b72d",
  1621 => x"831480f5",
  1622 => x"2d737081",
  1623 => x"055581b7",
  1624 => x"2d851480",
  1625 => x"f52d7370",
  1626 => x"81055581",
  1627 => x"b72d8714",
  1628 => x"80f52d73",
  1629 => x"70810555",
  1630 => x"81b72d89",
  1631 => x"1480f52d",
  1632 => x"73708105",
  1633 => x"5581b72d",
  1634 => x"8e1480f5",
  1635 => x"2d737081",
  1636 => x"055581b7",
  1637 => x"2d901480",
  1638 => x"f52d7370",
  1639 => x"81055581",
  1640 => x"b72d9214",
  1641 => x"80f52d73",
  1642 => x"70810555",
  1643 => x"81b72d94",
  1644 => x"1480f52d",
  1645 => x"73708105",
  1646 => x"5581b72d",
  1647 => x"961480f5",
  1648 => x"2d737081",
  1649 => x"055581b7",
  1650 => x"2d981480",
  1651 => x"f52d7370",
  1652 => x"81055581",
  1653 => x"b72d9c14",
  1654 => x"80f52d73",
  1655 => x"70810555",
  1656 => x"81b72d9e",
  1657 => x"1480f52d",
  1658 => x"7381b72d",
  1659 => x"7780d088",
  1660 => x"0c805372",
  1661 => x"80d1c40c",
  1662 => x"02a0050d",
  1663 => x"0402cc05",
  1664 => x"0d7e605e",
  1665 => x"5a800b80",
  1666 => x"d8e80880",
  1667 => x"d8ec0859",
  1668 => x"5c568058",
  1669 => x"80d8c808",
  1670 => x"782e81b8",
  1671 => x"38778f06",
  1672 => x"a0175754",
  1673 => x"73913880",
  1674 => x"d2b85276",
  1675 => x"51811757",
  1676 => x"a7ac2d80",
  1677 => x"d2b85680",
  1678 => x"7680f52d",
  1679 => x"56547474",
  1680 => x"2e833881",
  1681 => x"547481e5",
  1682 => x"2e80fd38",
  1683 => x"81707506",
  1684 => x"555c7380",
  1685 => x"2e80f138",
  1686 => x"8b1680f5",
  1687 => x"2d980659",
  1688 => x"7880e538",
  1689 => x"8b537c52",
  1690 => x"7551a8d0",
  1691 => x"2d80d1c4",
  1692 => x"0880d538",
  1693 => x"9c160851",
  1694 => x"b6f32d80",
  1695 => x"d1c40884",
  1696 => x"1b0c9a16",
  1697 => x"80e02d51",
  1698 => x"b7a42d80",
  1699 => x"d1c40880",
  1700 => x"d1c40888",
  1701 => x"1c0c80d1",
  1702 => x"c4085555",
  1703 => x"80d8c408",
  1704 => x"802e9938",
  1705 => x"941680e0",
  1706 => x"2d51b7a4",
  1707 => x"2d80d1c4",
  1708 => x"08902b83",
  1709 => x"fff00a06",
  1710 => x"70165154",
  1711 => x"73881b0c",
  1712 => x"787a0c7b",
  1713 => x"54b69004",
  1714 => x"81185880",
  1715 => x"d8c80878",
  1716 => x"26feca38",
  1717 => x"80d8c408",
  1718 => x"802eb338",
  1719 => x"7a51b0c9",
  1720 => x"2d80d1c4",
  1721 => x"0880d1c4",
  1722 => x"0880ffff",
  1723 => x"fff80655",
  1724 => x"5b7380ff",
  1725 => x"fffff82e",
  1726 => x"953880d1",
  1727 => x"c408fe05",
  1728 => x"80d8bc08",
  1729 => x"2980d8d0",
  1730 => x"080557b4",
  1731 => x"92048054",
  1732 => x"7380d1c4",
  1733 => x"0c02b405",
  1734 => x"0d0402f4",
  1735 => x"050d7470",
  1736 => x"08810571",
  1737 => x"0c700880",
  1738 => x"d8c00806",
  1739 => x"5353718f",
  1740 => x"38881308",
  1741 => x"51b0c92d",
  1742 => x"80d1c408",
  1743 => x"88140c81",
  1744 => x"0b80d1c4",
  1745 => x"0c028c05",
  1746 => x"0d0402f0",
  1747 => x"050d7588",
  1748 => x"1108fe05",
  1749 => x"80d8bc08",
  1750 => x"2980d8d0",
  1751 => x"08117208",
  1752 => x"80d8c008",
  1753 => x"06057955",
  1754 => x"535454a7",
  1755 => x"ac2d0290",
  1756 => x"050d0402",
  1757 => x"f4050d74",
  1758 => x"70882a83",
  1759 => x"fe800670",
  1760 => x"72982a07",
  1761 => x"72882b87",
  1762 => x"fc808006",
  1763 => x"73982b81",
  1764 => x"f00a0671",
  1765 => x"73070780",
  1766 => x"d1c40c56",
  1767 => x"51535102",
  1768 => x"8c050d04",
  1769 => x"02f8050d",
  1770 => x"028e0580",
  1771 => x"f52d7488",
  1772 => x"2b077083",
  1773 => x"ffff0680",
  1774 => x"d1c40c51",
  1775 => x"0288050d",
  1776 => x"0402f405",
  1777 => x"0d747678",
  1778 => x"53545280",
  1779 => x"71259738",
  1780 => x"72708105",
  1781 => x"5480f52d",
  1782 => x"72708105",
  1783 => x"5481b72d",
  1784 => x"ff115170",
  1785 => x"eb388072",
  1786 => x"81b72d02",
  1787 => x"8c050d04",
  1788 => x"02e8050d",
  1789 => x"77568070",
  1790 => x"56547376",
  1791 => x"24b63880",
  1792 => x"d8c80874",
  1793 => x"2eae3873",
  1794 => x"51b1c22d",
  1795 => x"80d1c408",
  1796 => x"80d1c408",
  1797 => x"09810570",
  1798 => x"80d1c408",
  1799 => x"079f2a77",
  1800 => x"05811757",
  1801 => x"57535374",
  1802 => x"76248938",
  1803 => x"80d8c808",
  1804 => x"7426d438",
  1805 => x"7280d1c4",
  1806 => x"0c029805",
  1807 => x"0d0402ec",
  1808 => x"050d80d1",
  1809 => x"c0081751",
  1810 => x"b7f02d80",
  1811 => x"d1c40855",
  1812 => x"80d1c408",
  1813 => x"802ea238",
  1814 => x"8b5380d1",
  1815 => x"c4085280",
  1816 => x"d6b851b7",
  1817 => x"c12d80d8",
  1818 => x"f4085473",
  1819 => x"802e8a38",
  1820 => x"88155280",
  1821 => x"d6b85173",
  1822 => x"2d029405",
  1823 => x"0d0402dc",
  1824 => x"050d8070",
  1825 => x"5a557480",
  1826 => x"d1c00825",
  1827 => x"b43880d8",
  1828 => x"c808752e",
  1829 => x"ac387851",
  1830 => x"b1c22d80",
  1831 => x"d1c40809",
  1832 => x"81057080",
  1833 => x"d1c40807",
  1834 => x"9f2a7605",
  1835 => x"811b5b56",
  1836 => x"547480d1",
  1837 => x"c0082589",
  1838 => x"3880d8c8",
  1839 => x"087926d6",
  1840 => x"38805578",
  1841 => x"80d8c808",
  1842 => x"2781db38",
  1843 => x"7851b1c2",
  1844 => x"2d80d1c4",
  1845 => x"08802e81",
  1846 => x"ad3880d1",
  1847 => x"c4088b05",
  1848 => x"80f52d70",
  1849 => x"842a7081",
  1850 => x"06771078",
  1851 => x"842b80d6",
  1852 => x"b80b80f5",
  1853 => x"2d5c5c53",
  1854 => x"51555673",
  1855 => x"802e80cb",
  1856 => x"38741682",
  1857 => x"2bbbca0b",
  1858 => x"80d09412",
  1859 => x"0c547775",
  1860 => x"311080d8",
  1861 => x"f8115556",
  1862 => x"90747081",
  1863 => x"055681b7",
  1864 => x"2da07481",
  1865 => x"b72d7681",
  1866 => x"ff068116",
  1867 => x"58547380",
  1868 => x"2e8a389c",
  1869 => x"5380d6b8",
  1870 => x"52bac304",
  1871 => x"8b5380d1",
  1872 => x"c4085280",
  1873 => x"d8fa1651",
  1874 => x"bafe0474",
  1875 => x"16822bb8",
  1876 => x"be0b80d0",
  1877 => x"94120c54",
  1878 => x"7681ff06",
  1879 => x"81165854",
  1880 => x"73802e8a",
  1881 => x"389c5380",
  1882 => x"d6b852ba",
  1883 => x"f5048b53",
  1884 => x"80d1c408",
  1885 => x"52777531",
  1886 => x"1080d8f8",
  1887 => x"05517655",
  1888 => x"b7c12dbb",
  1889 => x"9b047490",
  1890 => x"29753170",
  1891 => x"1080d8f8",
  1892 => x"05515480",
  1893 => x"d1c40874",
  1894 => x"81b72d81",
  1895 => x"1959748b",
  1896 => x"24a338b9",
  1897 => x"c3047490",
  1898 => x"29753170",
  1899 => x"1080d8f8",
  1900 => x"058c7731",
  1901 => x"57515480",
  1902 => x"7481b72d",
  1903 => x"9e14ff16",
  1904 => x"565474f3",
  1905 => x"3802a405",
  1906 => x"0d0402fc",
  1907 => x"050d80d1",
  1908 => x"c0081351",
  1909 => x"b7f02d80",
  1910 => x"d1c40880",
  1911 => x"2e893880",
  1912 => x"d1c40851",
  1913 => x"a98f2d80",
  1914 => x"0b80d1c0",
  1915 => x"0cb8fe2d",
  1916 => x"93e02d02",
  1917 => x"84050d04",
  1918 => x"02fc050d",
  1919 => x"725170fd",
  1920 => x"2eb03870",
  1921 => x"fd248a38",
  1922 => x"70fc2e80",
  1923 => x"cc38bce3",
  1924 => x"0470fe2e",
  1925 => x"b73870ff",
  1926 => x"2e098106",
  1927 => x"80c53880",
  1928 => x"d1c00851",
  1929 => x"70802ebb",
  1930 => x"38ff1180",
  1931 => x"d1c00cbc",
  1932 => x"e30480d1",
  1933 => x"c008f405",
  1934 => x"7080d1c0",
  1935 => x"0c517080",
  1936 => x"25a13880",
  1937 => x"0b80d1c0",
  1938 => x"0cbce304",
  1939 => x"80d1c008",
  1940 => x"810580d1",
  1941 => x"c00cbce3",
  1942 => x"0480d1c0",
  1943 => x"088c0580",
  1944 => x"d1c00cb8",
  1945 => x"fe2d93e0",
  1946 => x"2d028405",
  1947 => x"0d0402fc",
  1948 => x"050d800b",
  1949 => x"80d1c00c",
  1950 => x"b8fe2d92",
  1951 => x"ce2d80d1",
  1952 => x"c40880d1",
  1953 => x"b00c80d0",
  1954 => x"8c519586",
  1955 => x"2d028405",
  1956 => x"0d0402fc",
  1957 => x"050d810b",
  1958 => x"80c9800c",
  1959 => x"7251bcee",
  1960 => x"2d028405",
  1961 => x"0d0402fc",
  1962 => x"050d800b",
  1963 => x"80c9800c",
  1964 => x"7251bcee",
  1965 => x"2d028405",
  1966 => x"0d047180",
  1967 => x"d8f40c04",
  1968 => x"00ffffff",
  1969 => x"ff00ffff",
  1970 => x"ffff00ff",
  1971 => x"ffffff00",
  1972 => x"4b455953",
  1973 => x"50312020",
  1974 => x"20202000",
  1975 => x"00000000",
  1976 => x"4b455953",
  1977 => x"50322020",
  1978 => x"20202000",
  1979 => x"00000000",
  1980 => x"3d3d2056",
  1981 => x"6964656f",
  1982 => x"70616320",
  1983 => x"666f7220",
  1984 => x"5a58444f",
  1985 => x"53203d3d",
  1986 => x"00000000",
  1987 => x"3d3d3d3d",
  1988 => x"3d3d3d3d",
  1989 => x"3d3d3d3d",
  1990 => x"3d3d3d3d",
  1991 => x"3d3d3d3d",
  1992 => x"3d3d3d3d",
  1993 => x"00000000",
  1994 => x"52657365",
  1995 => x"74000000",
  1996 => x"5363616e",
  1997 => x"6c696e65",
  1998 => x"73000000",
  1999 => x"53776170",
  2000 => x"206a6f79",
  2001 => x"73746963",
  2002 => x"6b730000",
  2003 => x"4a6f696e",
  2004 => x"206a6f79",
  2005 => x"73746963",
  2006 => x"6b730000",
  2007 => x"4c6f6164",
  2008 => x"20636174",
  2009 => x"72696467",
  2010 => x"6520524f",
  2011 => x"4d201000",
  2012 => x"4c6f6164",
  2013 => x"20564443",
  2014 => x"20666f6e",
  2015 => x"74201000",
  2016 => x"48656c70",
  2017 => x"00000000",
  2018 => x"45786974",
  2019 => x"00000000",
  2020 => x"54686520",
  2021 => x"766f6963",
  2022 => x"653a204f",
  2023 => x"66660000",
  2024 => x"54686520",
  2025 => x"766f6963",
  2026 => x"653a204f",
  2027 => x"6e000000",
  2028 => x"436f6c6f",
  2029 => x"72206d6f",
  2030 => x"64653a20",
  2031 => x"436f6c6f",
  2032 => x"72000000",
  2033 => x"436f6c6f",
  2034 => x"72206d6f",
  2035 => x"64653a20",
  2036 => x"4d6f6e6f",
  2037 => x"6368726f",
  2038 => x"6d650000",
  2039 => x"436f6c6f",
  2040 => x"72206d6f",
  2041 => x"64653a20",
  2042 => x"47726565",
  2043 => x"6e207068",
  2044 => x"6f737068",
  2045 => x"6f720000",
  2046 => x"436f6c6f",
  2047 => x"72206d6f",
  2048 => x"64653a20",
  2049 => x"416d6265",
  2050 => x"72206d6f",
  2051 => x"6e6f6368",
  2052 => x"726f6d65",
  2053 => x"00000000",
  2054 => x"4d6f6465",
  2055 => x"3a204f64",
  2056 => x"79737365",
  2057 => x"79322028",
  2058 => x"4e545343",
  2059 => x"29000000",
  2060 => x"4d6f6465",
  2061 => x"3a205669",
  2062 => x"64656f70",
  2063 => x"61632028",
  2064 => x"50414c29",
  2065 => x"00000000",
  2066 => x"3d3d2056",
  2067 => x"6964656f",
  2068 => x"70616320",
  2069 => x"666f7220",
  2070 => x"5a58554e",
  2071 => x"4f203d3d",
  2072 => x"00000000",
  2073 => x"5a58554e",
  2074 => x"4f3a2073",
  2075 => x"696e676c",
  2076 => x"65206a6f",
  2077 => x"79737469",
  2078 => x"636b0000",
  2079 => x"5a58554e",
  2080 => x"4f3a2032",
  2081 => x"206a6f79",
  2082 => x"73746963",
  2083 => x"6b207370",
  2084 => x"6c697474",
  2085 => x"65720000",
  2086 => x"5a58554e",
  2087 => x"4f3a2032",
  2088 => x"206a6f79",
  2089 => x"73746963",
  2090 => x"6b205647",
  2091 => x"41324d00",
  2092 => x"524f4d20",
  2093 => x"6c6f6164",
  2094 => x"696e6720",
  2095 => x"6661696c",
  2096 => x"65640000",
  2097 => x"4f4b0000",
  2098 => x"3d3d3d20",
  2099 => x"56696465",
  2100 => x"6f706163",
  2101 => x"20537065",
  2102 => x"6369616c",
  2103 => x"2048454c",
  2104 => x"50203d3d",
  2105 => x"3d000000",
  2106 => x"3d3d3d3d",
  2107 => x"3d3d3d3d",
  2108 => x"3d3d3d3d",
  2109 => x"3d3d3d3d",
  2110 => x"3d3d3d3d",
  2111 => x"3d3d3d3d",
  2112 => x"3d3d3d3d",
  2113 => x"3d3d0000",
  2114 => x"5363726f",
  2115 => x"6c6c204c",
  2116 => x"6f636b3a",
  2117 => x"20636861",
  2118 => x"6e676520",
  2119 => x"62657477",
  2120 => x"65656e00",
  2121 => x"52474220",
  2122 => x"616e6420",
  2123 => x"56474120",
  2124 => x"76696465",
  2125 => x"6f206d6f",
  2126 => x"64650000",
  2127 => x"46333a20",
  2128 => x"536f6674",
  2129 => x"20526573",
  2130 => x"65740000",
  2131 => x"4374726c",
  2132 => x"2b416c74",
  2133 => x"2b426163",
  2134 => x"6b737061",
  2135 => x"63653a20",
  2136 => x"48617264",
  2137 => x"20726573",
  2138 => x"65740000",
  2139 => x"45736320",
  2140 => x"6f72206a",
  2141 => x"6f797374",
  2142 => x"69636b20",
  2143 => x"62742e32",
  2144 => x"3a20746f",
  2145 => x"2073686f",
  2146 => x"77000000",
  2147 => x"6f722068",
  2148 => x"69646520",
  2149 => x"74686520",
  2150 => x"6f707469",
  2151 => x"6f6e7320",
  2152 => x"6d656e75",
  2153 => x"2e000000",
  2154 => x"57415344",
  2155 => x"202f2063",
  2156 => x"7572736f",
  2157 => x"72206b65",
  2158 => x"7973202f",
  2159 => x"206a6f79",
  2160 => x"73746963",
  2161 => x"6b000000",
  2162 => x"746f2073",
  2163 => x"656c6563",
  2164 => x"74206d65",
  2165 => x"6e75206f",
  2166 => x"7074696f",
  2167 => x"6e2e0000",
  2168 => x"456e7465",
  2169 => x"72202f20",
  2170 => x"46697265",
  2171 => x"20746f20",
  2172 => x"63686f6f",
  2173 => x"7365206f",
  2174 => x"7074696f",
  2175 => x"6e2e0000",
  2176 => x"496e206d",
  2177 => x"6f737420",
  2178 => x"67616d65",
  2179 => x"73207072",
  2180 => x"65737320",
  2181 => x"302d3920",
  2182 => x"61667465",
  2183 => x"72000000",
  2184 => x"6c6f6164",
  2185 => x"696e6720",
  2186 => x"6120524f",
  2187 => x"4d20746f",
  2188 => x"20706c61",
  2189 => x"79207468",
  2190 => x"65206761",
  2191 => x"6d650000",
  2192 => x"3d3d3d20",
  2193 => x"56696465",
  2194 => x"6f706163",
  2195 => x"20436f72",
  2196 => x"65204372",
  2197 => x"65646974",
  2198 => x"73203d3d",
  2199 => x"3d000000",
  2200 => x"3d3d3d3d",
  2201 => x"3d3d3d3d",
  2202 => x"3d3d3d3d",
  2203 => x"3d3d3d3d",
  2204 => x"3d3d3d3d",
  2205 => x"3d3d3d3d",
  2206 => x"3d3d3d3d",
  2207 => x"3d000000",
  2208 => x"5068696c",
  2209 => x"69707320",
  2210 => x"56696465",
  2211 => x"6f706163",
  2212 => x"202f204d",
  2213 => x"61676e61",
  2214 => x"766f7800",
  2215 => x"4f647973",
  2216 => x"73657932",
  2217 => x"20636f72",
  2218 => x"6520666f",
  2219 => x"72205a58",
  2220 => x"554e4f2c",
  2221 => x"205a5844",
  2222 => x"4f530000",
  2223 => x"616e6420",
  2224 => x"5a58444f",
  2225 => x"532b2062",
  2226 => x"6f617264",
  2227 => x"732e0000",
  2228 => x"4f726967",
  2229 => x"696e616c",
  2230 => x"20636f72",
  2231 => x"65206279",
  2232 => x"3a41726e",
  2233 => x"696d204c",
  2234 => x"61657567",
  2235 => x"65720000",
  2236 => x"506f7274",
  2237 => x"206d6164",
  2238 => x"65206279",
  2239 => x"3a20796f",
  2240 => x"6d626f70",
  2241 => x"72696d65",
  2242 => x"2c200000",
  2243 => x"2072616d",
  2244 => x"70613036",
  2245 => x"392c206e",
  2246 => x"6575726f",
  2247 => x"72756c65",
  2248 => x"7a2c2041",
  2249 => x"6e746f6e",
  2250 => x"696f0000",
  2251 => x"2053616e",
  2252 => x"6368657a",
  2253 => x"2c204176",
  2254 => x"6c697841",
  2255 => x"2c204d65",
  2256 => x"6a696173",
  2257 => x"33442c20",
  2258 => x"00000000",
  2259 => x"2057696c",
  2260 => x"636f3230",
  2261 => x"30392061",
  2262 => x"6e642042",
  2263 => x"656e6974",
  2264 => x"6f737300",
  2265 => x"53706563",
  2266 => x"69616c20",
  2267 => x"5468616e",
  2268 => x"6b732074",
  2269 => x"6f3a2052",
  2270 => x"656e6520",
  2271 => x"76616e20",
  2272 => x"00000000",
  2273 => x"2064656e",
  2274 => x"20456e64",
  2275 => x"656e2066",
  2276 => x"6f722068",
  2277 => x"69732069",
  2278 => x"6e666f20",
  2279 => x"6f6e2000",
  2280 => x"20766964",
  2281 => x"656f7061",
  2282 => x"632e6e6c",
  2283 => x"00000000",
  2284 => x"496e6974",
  2285 => x"69616c69",
  2286 => x"7a696e67",
  2287 => x"20534420",
  2288 => x"63617264",
  2289 => x"0a000000",
  2290 => x"16200000",
  2291 => x"14200000",
  2292 => x"15200000",
  2293 => x"53442069",
  2294 => x"6e69742e",
  2295 => x"2e2e0a00",
  2296 => x"53442063",
  2297 => x"61726420",
  2298 => x"72657365",
  2299 => x"74206661",
  2300 => x"696c6564",
  2301 => x"210a0000",
  2302 => x"53444843",
  2303 => x"20657272",
  2304 => x"6f72210a",
  2305 => x"00000000",
  2306 => x"57726974",
  2307 => x"65206661",
  2308 => x"696c6564",
  2309 => x"0a000000",
  2310 => x"52656164",
  2311 => x"20666169",
  2312 => x"6c65640a",
  2313 => x"00000000",
  2314 => x"43617264",
  2315 => x"20696e69",
  2316 => x"74206661",
  2317 => x"696c6564",
  2318 => x"0a000000",
  2319 => x"46415431",
  2320 => x"36202020",
  2321 => x"00000000",
  2322 => x"46415433",
  2323 => x"32202020",
  2324 => x"00000000",
  2325 => x"4e6f2070",
  2326 => x"61727469",
  2327 => x"74696f6e",
  2328 => x"20736967",
  2329 => x"0a000000",
  2330 => x"42616420",
  2331 => x"70617274",
  2332 => x"0a000000",
  2333 => x"4261636b",
  2334 => x"00000000",
  2335 => x"00000002",
  2336 => x"00000000",
  2337 => x"00000010",
  2338 => x"00000002",
  2339 => x"00001ef0",
  2340 => x"000003ab",
  2341 => x"00000002",
  2342 => x"00001f0c",
  2343 => x"000003ab",
  2344 => x"00000002",
  2345 => x"00001f28",
  2346 => x"0000037f",
  2347 => x"00000001",
  2348 => x"00001f30",
  2349 => x"00000000",
  2350 => x"00000001",
  2351 => x"00001f3c",
  2352 => x"00000001",
  2353 => x"00000001",
  2354 => x"00001f4c",
  2355 => x"00000002",
  2356 => x"00000002",
  2357 => x"00001f5c",
  2358 => x"00001ea6",
  2359 => x"00000002",
  2360 => x"00001f70",
  2361 => x"00001e92",
  2362 => x"00000003",
  2363 => x"00002548",
  2364 => x"00000002",
  2365 => x"00000003",
  2366 => x"00002538",
  2367 => x"00000004",
  2368 => x"00000003",
  2369 => x"00002530",
  2370 => x"00000002",
  2371 => x"00000002",
  2372 => x"00001f80",
  2373 => x"000003c6",
  2374 => x"00000002",
  2375 => x"00001f88",
  2376 => x"0000096b",
  2377 => x"00000000",
  2378 => x"00000000",
  2379 => x"00000000",
  2380 => x"00001f90",
  2381 => x"00001fa0",
  2382 => x"00001fb0",
  2383 => x"00001fc4",
  2384 => x"00001fdc",
  2385 => x"00001ff8",
  2386 => x"00002018",
  2387 => x"00002030",
  2388 => x"00000002",
  2389 => x"00002048",
  2390 => x"000003ab",
  2391 => x"00000002",
  2392 => x"00001f0c",
  2393 => x"000003ab",
  2394 => x"00000002",
  2395 => x"00001f28",
  2396 => x"0000037f",
  2397 => x"00000001",
  2398 => x"00001f30",
  2399 => x"00000000",
  2400 => x"00000001",
  2401 => x"00001f3c",
  2402 => x"00000001",
  2403 => x"00000001",
  2404 => x"00001f4c",
  2405 => x"00000002",
  2406 => x"00000002",
  2407 => x"00001f5c",
  2408 => x"00001ea6",
  2409 => x"00000002",
  2410 => x"00001f70",
  2411 => x"00001e92",
  2412 => x"00000003",
  2413 => x"00002548",
  2414 => x"00000002",
  2415 => x"00000003",
  2416 => x"00002538",
  2417 => x"00000004",
  2418 => x"00000003",
  2419 => x"000025f8",
  2420 => x"00000003",
  2421 => x"00000002",
  2422 => x"00001f80",
  2423 => x"000003c6",
  2424 => x"00000002",
  2425 => x"00001f88",
  2426 => x"0000096b",
  2427 => x"00000000",
  2428 => x"00000000",
  2429 => x"00000000",
  2430 => x"00002064",
  2431 => x"0000207c",
  2432 => x"00002098",
  2433 => x"00000004",
  2434 => x"000020b0",
  2435 => x"00002604",
  2436 => x"00000004",
  2437 => x"000020c4",
  2438 => x"000028ec",
  2439 => x"00000000",
  2440 => x"00000000",
  2441 => x"00000000",
  2442 => x"00000002",
  2443 => x"000020c8",
  2444 => x"000003aa",
  2445 => x"00000002",
  2446 => x"000020e8",
  2447 => x"000003aa",
  2448 => x"00000002",
  2449 => x"00002108",
  2450 => x"000003aa",
  2451 => x"00000002",
  2452 => x"00002124",
  2453 => x"000003aa",
  2454 => x"00000002",
  2455 => x"0000213c",
  2456 => x"000003aa",
  2457 => x"00000002",
  2458 => x"0000214c",
  2459 => x"000003aa",
  2460 => x"00000002",
  2461 => x"0000216c",
  2462 => x"000003aa",
  2463 => x"00000002",
  2464 => x"0000218c",
  2465 => x"000003aa",
  2466 => x"00000002",
  2467 => x"000021a8",
  2468 => x"000003aa",
  2469 => x"00000002",
  2470 => x"000021c8",
  2471 => x"000003aa",
  2472 => x"00000002",
  2473 => x"000021e0",
  2474 => x"000003aa",
  2475 => x"00000002",
  2476 => x"00002200",
  2477 => x"000003aa",
  2478 => x"00000002",
  2479 => x"00002220",
  2480 => x"000003aa",
  2481 => x"00000004",
  2482 => x"000020c4",
  2483 => x"000028ec",
  2484 => x"00000000",
  2485 => x"00000000",
  2486 => x"00000000",
  2487 => x"00000002",
  2488 => x"00002240",
  2489 => x"000003aa",
  2490 => x"00000002",
  2491 => x"00002260",
  2492 => x"000003aa",
  2493 => x"00000002",
  2494 => x"00002280",
  2495 => x"000003aa",
  2496 => x"00000002",
  2497 => x"0000229c",
  2498 => x"000003aa",
  2499 => x"00000002",
  2500 => x"000022bc",
  2501 => x"000003aa",
  2502 => x"00000002",
  2503 => x"000022d0",
  2504 => x"000003aa",
  2505 => x"00000002",
  2506 => x"000022f0",
  2507 => x"000003aa",
  2508 => x"00000002",
  2509 => x"0000230c",
  2510 => x"000003aa",
  2511 => x"00000002",
  2512 => x"0000232c",
  2513 => x"000003aa",
  2514 => x"00000002",
  2515 => x"0000234c",
  2516 => x"000003aa",
  2517 => x"00000002",
  2518 => x"00002364",
  2519 => x"000003aa",
  2520 => x"00000002",
  2521 => x"00002384",
  2522 => x"000003aa",
  2523 => x"00000002",
  2524 => x"000023a0",
  2525 => x"000003aa",
  2526 => x"00000004",
  2527 => x"000020c4",
  2528 => x"000028ec",
  2529 => x"00000000",
  2530 => x"00000000",
  2531 => x"00000000",
  2532 => x"00000000",
  2533 => x"00000000",
  2534 => x"00000000",
  2535 => x"00000000",
  2536 => x"00000000",
  2537 => x"00000000",
  2538 => x"00000000",
  2539 => x"00000000",
  2540 => x"00000000",
  2541 => x"00000000",
  2542 => x"00000000",
  2543 => x"00000000",
  2544 => x"00000000",
  2545 => x"00000000",
  2546 => x"00000000",
  2547 => x"00000000",
  2548 => x"00000000",
  2549 => x"00000000",
  2550 => x"00000006",
  2551 => x"00000043",
  2552 => x"00000042",
  2553 => x"0000003b",
  2554 => x"0000004b",
  2555 => x"00000033",
  2556 => x"0000001d",
  2557 => x"0000001b",
  2558 => x"0000001c",
  2559 => x"00000023",
  2560 => x"0000002b",
  2561 => x"00000000",
  2562 => x"00000000",
  2563 => x"00000002",
  2564 => x"00002c78",
  2565 => x"00001c3e",
  2566 => x"00000002",
  2567 => x"00002c96",
  2568 => x"00001c3e",
  2569 => x"00000002",
  2570 => x"00002cb4",
  2571 => x"00001c3e",
  2572 => x"00000002",
  2573 => x"00002cd2",
  2574 => x"00001c3e",
  2575 => x"00000002",
  2576 => x"00002cf0",
  2577 => x"00001c3e",
  2578 => x"00000002",
  2579 => x"00002d0e",
  2580 => x"00001c3e",
  2581 => x"00000002",
  2582 => x"00002d2c",
  2583 => x"00001c3e",
  2584 => x"00000002",
  2585 => x"00002d4a",
  2586 => x"00001c3e",
  2587 => x"00000002",
  2588 => x"00002d68",
  2589 => x"00001c3e",
  2590 => x"00000002",
  2591 => x"00002d86",
  2592 => x"00001c3e",
  2593 => x"00000002",
  2594 => x"00002da4",
  2595 => x"00001c3e",
  2596 => x"00000002",
  2597 => x"00002dc2",
  2598 => x"00001c3e",
  2599 => x"00000002",
  2600 => x"00002de0",
  2601 => x"00001c3e",
  2602 => x"00000004",
  2603 => x"00002474",
  2604 => x"00000000",
  2605 => x"00000000",
  2606 => x"00000000",
  2607 => x"00001df8",
  2608 => x"00000000",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memAWriteEnable = '1') and (from_zpu.memBWriteEnable = '1') and (from_zpu.memAAddr=from_zpu.memBAddr) and (from_zpu.memAWrite/=from_zpu.memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (from_zpu.memAWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memAWrite;
			to_zpu.memARead <= from_zpu.memAWrite;
		else
			to_zpu.memARead <= ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memBWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memBWrite;
			to_zpu.memBRead <= from_zpu.memBWrite;
		else
			to_zpu.memBRead <= ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;


end arch;

