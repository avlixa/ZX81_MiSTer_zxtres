-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Alastair M. Robinson for the ZPUFlex project.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.zpupkg.all;

entity CtrlROM_ROM is
generic
	(
		maxAddrBitBRAM : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_zpu : in ZPU_ToROM;
	to_zpu : out ZPU_FromROM
);
end CtrlROM_ROM;

architecture arch of CtrlROM_ROM is

type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"0b0b0b0b",
     1 => x"8c0b0b0b",
     2 => x"0b81e004",
     3 => x"0b0b0b0b",
     4 => x"8c04ff0d",
     5 => x"80040400",
     6 => x"00000016",
     7 => x"00000000",
     8 => x"0b0b80d2",
     9 => x"bc080b0b",
    10 => x"80d2c008",
    11 => x"0b0b80d2",
    12 => x"c4080b0b",
    13 => x"0b0b9808",
    14 => x"2d0b0b80",
    15 => x"d2c40c0b",
    16 => x"0b80d2c0",
    17 => x"0c0b0b80",
    18 => x"d2bc0c04",
    19 => x"00000000",
    20 => x"00000000",
    21 => x"00000000",
    22 => x"00000000",
    23 => x"00000000",
    24 => x"71fd0608",
    25 => x"72830609",
    26 => x"81058205",
    27 => x"832b2a83",
    28 => x"ffff0652",
    29 => x"0471fc06",
    30 => x"08728306",
    31 => x"09810583",
    32 => x"05101010",
    33 => x"2a81ff06",
    34 => x"520471fd",
    35 => x"060883ff",
    36 => x"ff738306",
    37 => x"09810582",
    38 => x"05832b2b",
    39 => x"09067383",
    40 => x"ffff0673",
    41 => x"83060981",
    42 => x"05820583",
    43 => x"2b0b2b07",
    44 => x"72fc060c",
    45 => x"51510471",
    46 => x"fc06080b",
    47 => x"0b0bbd88",
    48 => x"73830610",
    49 => x"10050806",
    50 => x"7381ff06",
    51 => x"73830609",
    52 => x"81058305",
    53 => x"1010102b",
    54 => x"0772fc06",
    55 => x"0c515104",
    56 => x"80d2bc70",
    57 => x"80dcfc27",
    58 => x"8b388071",
    59 => x"70840553",
    60 => x"0c81e304",
    61 => x"8c518a91",
    62 => x"0402fc05",
    63 => x"0df88051",
    64 => x"8f0b80d2",
    65 => x"cc0c9f0b",
    66 => x"80d2d00c",
    67 => x"a0717081",
    68 => x"05533480",
    69 => x"d2d008ff",
    70 => x"0580d2d0",
    71 => x"0c80d2d0",
    72 => x"088025e8",
    73 => x"3880d2cc",
    74 => x"08ff0580",
    75 => x"d2cc0c80",
    76 => x"d2cc0880",
    77 => x"25d03880",
    78 => x"0b80d2d0",
    79 => x"0c800b80",
    80 => x"d2cc0c02",
    81 => x"84050d04",
    82 => x"02f0050d",
    83 => x"f88053f8",
    84 => x"a05483bf",
    85 => x"52737081",
    86 => x"05553351",
    87 => x"70737081",
    88 => x"055534ff",
    89 => x"12527180",
    90 => x"25eb38fb",
    91 => x"c0539f52",
    92 => x"a0737081",
    93 => x"055534ff",
    94 => x"12527180",
    95 => x"25f23802",
    96 => x"90050d04",
    97 => x"02f4050d",
    98 => x"74538e0b",
    99 => x"80d2cc08",
   100 => x"25913882",
   101 => x"c82d80d2",
   102 => x"cc08ff05",
   103 => x"80d2cc0c",
   104 => x"838a0480",
   105 => x"d2cc0880",
   106 => x"d2d00853",
   107 => x"51728a2e",
   108 => x"098106be",
   109 => x"38715171",
   110 => x"9f24a438",
   111 => x"80d2cc08",
   112 => x"a02911f8",
   113 => x"80115151",
   114 => x"a0713480",
   115 => x"d2d00881",
   116 => x"0580d2d0",
   117 => x"0c80d2d0",
   118 => x"08519f71",
   119 => x"25de3880",
   120 => x"0b80d2d0",
   121 => x"0c80d2cc",
   122 => x"08810580",
   123 => x"d2cc0c84",
   124 => x"880470a0",
   125 => x"2912f880",
   126 => x"11515172",
   127 => x"713480d2",
   128 => x"d0088105",
   129 => x"80d2d00c",
   130 => x"80d2d008",
   131 => x"a02e0981",
   132 => x"06913880",
   133 => x"0b80d2d0",
   134 => x"0c80d2cc",
   135 => x"08810580",
   136 => x"d2cc0c02",
   137 => x"8c050d04",
   138 => x"02f4050d",
   139 => x"74537270",
   140 => x"81055433",
   141 => x"5271802e",
   142 => x"89387151",
   143 => x"83842d84",
   144 => x"ae04810b",
   145 => x"80d2bc0c",
   146 => x"028c050d",
   147 => x"0402e805",
   148 => x"0d777956",
   149 => x"56880bfc",
   150 => x"1677712c",
   151 => x"8f065452",
   152 => x"54805372",
   153 => x"72259538",
   154 => x"7153fbe0",
   155 => x"14518771",
   156 => x"348114ff",
   157 => x"14545472",
   158 => x"f1387153",
   159 => x"f9157671",
   160 => x"2c870653",
   161 => x"5171802e",
   162 => x"8b38fbe0",
   163 => x"14517171",
   164 => x"34811454",
   165 => x"728e2495",
   166 => x"388f7331",
   167 => x"53fbe014",
   168 => x"51a07134",
   169 => x"8114ff14",
   170 => x"545472f1",
   171 => x"38029805",
   172 => x"0d0402ec",
   173 => x"050d800b",
   174 => x"80d2d40c",
   175 => x"f68c08f6",
   176 => x"90087188",
   177 => x"2c565381",
   178 => x"ff065373",
   179 => x"73258938",
   180 => x"7254820b",
   181 => x"80d2d40c",
   182 => x"71882c72",
   183 => x"81ff0653",
   184 => x"55747225",
   185 => x"8d387180",
   186 => x"d2d40884",
   187 => x"0780d2d4",
   188 => x"0c557384",
   189 => x"2b75832b",
   190 => x"565483f4",
   191 => x"74258f38",
   192 => x"830b0b0b",
   193 => x"80c9dc0c",
   194 => x"818c5386",
   195 => x"9904810b",
   196 => x"0b0b80c9",
   197 => x"dc0c80c6",
   198 => x"530b0b80",
   199 => x"c9dc0881",
   200 => x"712bff05",
   201 => x"f6880cfc",
   202 => x"08757531",
   203 => x"ffb005ff",
   204 => x"1371712c",
   205 => x"ff941a70",
   206 => x"9f2a1170",
   207 => x"812c80d2",
   208 => x"d4085254",
   209 => x"51535753",
   210 => x"51525276",
   211 => x"802e8538",
   212 => x"70810751",
   213 => x"70f6940c",
   214 => x"72098105",
   215 => x"f6800c71",
   216 => x"098105f6",
   217 => x"840c0294",
   218 => x"050d0404",
   219 => x"02fc050d",
   220 => x"80cee051",
   221 => x"94b42d02",
   222 => x"84050d04",
   223 => x"02fc050d",
   224 => x"80c9e051",
   225 => x"94b42d02",
   226 => x"84050d04",
   227 => x"02fc050d",
   228 => x"80cdb851",
   229 => x"94b42d02",
   230 => x"84050d04",
   231 => x"02fc050d",
   232 => x"81808051",
   233 => x"c0115170",
   234 => x"fb380284",
   235 => x"050d0471",
   236 => x"812e0981",
   237 => x"06893881",
   238 => x"c30bec0c",
   239 => x"87c30483",
   240 => x"0bec0c87",
   241 => x"9c2d820b",
   242 => x"ec0c0491",
   243 => x"fc2d80d2",
   244 => x"bc0880cd",
   245 => x"a80c91fc",
   246 => x"2d80d2bc",
   247 => x"0880ccd4",
   248 => x"0c91fc2d",
   249 => x"80d2bc08",
   250 => x"80cff80c",
   251 => x"91fc2d80",
   252 => x"d2bc0880",
   253 => x"ced00c91",
   254 => x"fc2d80d2",
   255 => x"bc0880cb",
   256 => x"840c0402",
   257 => x"fc050d84",
   258 => x"bf51879c",
   259 => x"2dff1151",
   260 => x"708025f6",
   261 => x"38028405",
   262 => x"0d0402dc",
   263 => x"050d8059",
   264 => x"81840bec",
   265 => x"0c7a5280",
   266 => x"d2d851b3",
   267 => x"8c2d80d2",
   268 => x"bc08792e",
   269 => x"819b3880",
   270 => x"d2dc0854",
   271 => x"73852e09",
   272 => x"81068a38",
   273 => x"840bec0c",
   274 => x"815389d9",
   275 => x"0473f80c",
   276 => x"81a40bec",
   277 => x"0c88832d",
   278 => x"78ff1556",
   279 => x"5874802e",
   280 => x"8b388118",
   281 => x"75812a56",
   282 => x"5888dd04",
   283 => x"f7185881",
   284 => x"59807425",
   285 => x"80d738a4",
   286 => x"0bec0c77",
   287 => x"52745184",
   288 => x"cd2d80d3",
   289 => x"b45280d2",
   290 => x"d851b5ff",
   291 => x"2d80d2bc",
   292 => x"08802ea0",
   293 => x"3880d3b4",
   294 => x"5783fc56",
   295 => x"76708405",
   296 => x"5808e80c",
   297 => x"fc165675",
   298 => x"8025f138",
   299 => x"81a40bec",
   300 => x"0c89bc04",
   301 => x"80d2bc08",
   302 => x"59848054",
   303 => x"80d2d851",
   304 => x"b5cf2dfc",
   305 => x"80148116",
   306 => x"565488f1",
   307 => x"04840bec",
   308 => x"0c80d2dc",
   309 => x"08f80c78",
   310 => x"537280d2",
   311 => x"bc0c02a4",
   312 => x"050d0402",
   313 => x"f8050d73",
   314 => x"51889a2d",
   315 => x"80d2bc08",
   316 => x"5280d2bc",
   317 => x"08802e88",
   318 => x"3880cce4",
   319 => x"518a8404",
   320 => x"80ccc051",
   321 => x"94b42d71",
   322 => x"80d2bc0c",
   323 => x"0288050d",
   324 => x"0402f005",
   325 => x"0d800b80",
   326 => x"d2e40c88",
   327 => x"832d8151",
   328 => x"87af2d88",
   329 => x"832d8051",
   330 => x"87af2d88",
   331 => x"832d840b",
   332 => x"ec0c91cc",
   333 => x"2d8df72d",
   334 => x"81f92d83",
   335 => x"5291af2d",
   336 => x"815185b2",
   337 => x"2dff1252",
   338 => x"718025f1",
   339 => x"3880c40b",
   340 => x"ec0c80c7",
   341 => x"d45184a8",
   342 => x"2da9c42d",
   343 => x"80d2bc08",
   344 => x"802e82fc",
   345 => x"3881840b",
   346 => x"ec0c80d2",
   347 => x"e408bfff",
   348 => x"ff068780",
   349 => x"077080d2",
   350 => x"e40cfc0c",
   351 => x"80c7ec51",
   352 => x"889a2d80",
   353 => x"d2bc0880",
   354 => x"2e9d3880",
   355 => x"c7f85188",
   356 => x"9a2d80d2",
   357 => x"bc08802e",
   358 => x"8e3880c8",
   359 => x"8451889a",
   360 => x"2d80d2bc",
   361 => x"08883880",
   362 => x"c8905184",
   363 => x"a82d8051",
   364 => x"87af2d80",
   365 => x"5185b22d",
   366 => x"840bec0c",
   367 => x"89e351bc",
   368 => x"ff2d80d2",
   369 => x"e40880d0",
   370 => x"d00c80d2",
   371 => x"e408fc0c",
   372 => x"80cbd40b",
   373 => x"80d2e80c",
   374 => x"80cbd451",
   375 => x"94b42d80",
   376 => x"5187cb2d",
   377 => x"850b80d3",
   378 => x"a80c9285",
   379 => x"2d805185",
   380 => x"b22d9299",
   381 => x"2d8e832d",
   382 => x"94c72d80",
   383 => x"ca800b80",
   384 => x"f52d80ca",
   385 => x"8c0b80f5",
   386 => x"2d718a2b",
   387 => x"718b2b07",
   388 => x"80caa40b",
   389 => x"80f52d70",
   390 => x"8d2b7207",
   391 => x"80cabc0b",
   392 => x"80f52d70",
   393 => x"8e2b7207",
   394 => x"80caec0b",
   395 => x"80f52d70",
   396 => x"912b7207",
   397 => x"7080d2e4",
   398 => x"0c80d0d0",
   399 => x"08708106",
   400 => x"54525354",
   401 => x"52545253",
   402 => x"54555371",
   403 => x"802e8838",
   404 => x"73810780",
   405 => x"d2e40c72",
   406 => x"812a7081",
   407 => x"06515271",
   408 => x"802e8b38",
   409 => x"80d2e408",
   410 => x"820780d2",
   411 => x"e40c7282",
   412 => x"2a708106",
   413 => x"51527180",
   414 => x"2e8b3880",
   415 => x"d2e40884",
   416 => x"0780d2e4",
   417 => x"0c72832a",
   418 => x"70810651",
   419 => x"5271802e",
   420 => x"8b3880d2",
   421 => x"e4088807",
   422 => x"80d2e40c",
   423 => x"72842a70",
   424 => x"81065152",
   425 => x"71802e8b",
   426 => x"3880d2e4",
   427 => x"08900780",
   428 => x"d2e40c72",
   429 => x"852a7081",
   430 => x"06515271",
   431 => x"802e8b38",
   432 => x"80d2e408",
   433 => x"a00780d2",
   434 => x"e40c80d2",
   435 => x"e408fc0c",
   436 => x"865280d2",
   437 => x"bc088338",
   438 => x"845271ec",
   439 => x"0c8bf504",
   440 => x"800b80d2",
   441 => x"bc0c0290",
   442 => x"050d0471",
   443 => x"980c04ff",
   444 => x"b00880d2",
   445 => x"bc0c0481",
   446 => x"0bffb00c",
   447 => x"04800bff",
   448 => x"b00c0402",
   449 => x"f4050d8f",
   450 => x"910480d2",
   451 => x"bc0881f0",
   452 => x"2e098106",
   453 => x"8a38810b",
   454 => x"80d0c80c",
   455 => x"8f910480",
   456 => x"d2bc0881",
   457 => x"e02e0981",
   458 => x"068a3881",
   459 => x"0b80d0cc",
   460 => x"0c8f9104",
   461 => x"80d2bc08",
   462 => x"5280d0cc",
   463 => x"08802e89",
   464 => x"3880d2bc",
   465 => x"08818005",
   466 => x"5271842c",
   467 => x"728f0653",
   468 => x"5380d0c8",
   469 => x"08802e9a",
   470 => x"38728429",
   471 => x"80d08805",
   472 => x"72138171",
   473 => x"2b700973",
   474 => x"0806730c",
   475 => x"5153538f",
   476 => x"85047284",
   477 => x"2980d088",
   478 => x"05721383",
   479 => x"712b7208",
   480 => x"07720c53",
   481 => x"53800b80",
   482 => x"d0cc0c80",
   483 => x"0b80d0c8",
   484 => x"0c80d2ec",
   485 => x"5190982d",
   486 => x"80d2bc08",
   487 => x"ff24feea",
   488 => x"38800b80",
   489 => x"d2bc0c02",
   490 => x"8c050d04",
   491 => x"02f8050d",
   492 => x"80d08852",
   493 => x"8f518072",
   494 => x"70840554",
   495 => x"0cff1151",
   496 => x"708025f2",
   497 => x"38028805",
   498 => x"0d0402f0",
   499 => x"050d7551",
   500 => x"8dfd2d70",
   501 => x"822cfc06",
   502 => x"80d08811",
   503 => x"72109e06",
   504 => x"71087072",
   505 => x"2a708306",
   506 => x"82742b70",
   507 => x"09740676",
   508 => x"0c545156",
   509 => x"57535153",
   510 => x"8df72d71",
   511 => x"80d2bc0c",
   512 => x"0290050d",
   513 => x"0402fc05",
   514 => x"0d725180",
   515 => x"710c800b",
   516 => x"84120c02",
   517 => x"84050d04",
   518 => x"02f0050d",
   519 => x"75700884",
   520 => x"12085353",
   521 => x"53ff5471",
   522 => x"712ea838",
   523 => x"8dfd2d84",
   524 => x"13087084",
   525 => x"29148811",
   526 => x"70087081",
   527 => x"ff068418",
   528 => x"08811187",
   529 => x"06841a0c",
   530 => x"53515551",
   531 => x"51518df7",
   532 => x"2d715473",
   533 => x"80d2bc0c",
   534 => x"0290050d",
   535 => x"0402f405",
   536 => x"0d8dfd2d",
   537 => x"e008708b",
   538 => x"2a708106",
   539 => x"51525370",
   540 => x"802ea138",
   541 => x"80d2ec08",
   542 => x"70842980",
   543 => x"d2f40574",
   544 => x"81ff0671",
   545 => x"0c515180",
   546 => x"d2ec0881",
   547 => x"11870680",
   548 => x"d2ec0c51",
   549 => x"728c2c83",
   550 => x"ff0680d3",
   551 => x"940c800b",
   552 => x"80d3980c",
   553 => x"8def2d8d",
   554 => x"f72d028c",
   555 => x"050d0402",
   556 => x"fc050d8d",
   557 => x"fd2d810b",
   558 => x"80d3980c",
   559 => x"8df72d80",
   560 => x"d3980851",
   561 => x"70f93802",
   562 => x"84050d04",
   563 => x"02fc050d",
   564 => x"80d2ec51",
   565 => x"90852d8f",
   566 => x"ac2d90dd",
   567 => x"518deb2d",
   568 => x"0284050d",
   569 => x"0402fc05",
   570 => x"0d8fcf51",
   571 => x"879c2dff",
   572 => x"11517080",
   573 => x"25f63802",
   574 => x"84050d04",
   575 => x"80d3a008",
   576 => x"80d2bc0c",
   577 => x"0402fc05",
   578 => x"0d810b80",
   579 => x"d0fc0c81",
   580 => x"5185b22d",
   581 => x"0284050d",
   582 => x"0402fc05",
   583 => x"0d92a304",
   584 => x"8e832d80",
   585 => x"f6518fca",
   586 => x"2d80d2bc",
   587 => x"08f23880",
   588 => x"da518fca",
   589 => x"2d80d2bc",
   590 => x"08e63880",
   591 => x"d0f80851",
   592 => x"8fca2d80",
   593 => x"d2bc08d8",
   594 => x"3880d2bc",
   595 => x"0880d0fc",
   596 => x"0c80d2bc",
   597 => x"085185b2",
   598 => x"2d028405",
   599 => x"0d0402ec",
   600 => x"050d7654",
   601 => x"8052870b",
   602 => x"881580f5",
   603 => x"2d565374",
   604 => x"72248338",
   605 => x"a0537251",
   606 => x"83842d81",
   607 => x"128b1580",
   608 => x"f52d5452",
   609 => x"727225de",
   610 => x"38029405",
   611 => x"0d0402f0",
   612 => x"050d80d3",
   613 => x"a0085481",
   614 => x"f92d800b",
   615 => x"80d3a40c",
   616 => x"7308802e",
   617 => x"81893882",
   618 => x"0b80d2d0",
   619 => x"0c80d3a4",
   620 => x"088f0680",
   621 => x"d2cc0c73",
   622 => x"08527183",
   623 => x"2e963871",
   624 => x"83268938",
   625 => x"71812eb0",
   626 => x"38949804",
   627 => x"71852ea0",
   628 => x"38949804",
   629 => x"881480f5",
   630 => x"2d841508",
   631 => x"80c8a853",
   632 => x"545284a8",
   633 => x"2d718429",
   634 => x"13700852",
   635 => x"52949c04",
   636 => x"735192de",
   637 => x"2d949804",
   638 => x"80d0d008",
   639 => x"8815082c",
   640 => x"70810651",
   641 => x"5271802e",
   642 => x"883880c8",
   643 => x"ac519495",
   644 => x"0480c8b0",
   645 => x"5184a82d",
   646 => x"84140851",
   647 => x"84a82d80",
   648 => x"d3a40881",
   649 => x"0580d3a4",
   650 => x"0c8c1454",
   651 => x"93a00402",
   652 => x"90050d04",
   653 => x"7180d3a0",
   654 => x"0c938e2d",
   655 => x"80d3a408",
   656 => x"ff0580d3",
   657 => x"a80c0402",
   658 => x"e8050d80",
   659 => x"d3a00880",
   660 => x"d3ac0857",
   661 => x"5580f651",
   662 => x"8fca2d80",
   663 => x"d2bc0881",
   664 => x"2a708106",
   665 => x"51527180",
   666 => x"2ea23894",
   667 => x"f1048e83",
   668 => x"2d80f651",
   669 => x"8fca2d80",
   670 => x"d2bc08f2",
   671 => x"3880d0fc",
   672 => x"08813270",
   673 => x"80d0fc0c",
   674 => x"5185b22d",
   675 => x"800b80d3",
   676 => x"9c0c8c51",
   677 => x"8fca2d80",
   678 => x"d2bc0881",
   679 => x"2a708106",
   680 => x"51527180",
   681 => x"2e80d138",
   682 => x"80d0d408",
   683 => x"80d0e808",
   684 => x"80d0d40c",
   685 => x"80d0e80c",
   686 => x"80d0d808",
   687 => x"80d0ec08",
   688 => x"80d0d80c",
   689 => x"80d0ec0c",
   690 => x"80d0dc08",
   691 => x"80d0f008",
   692 => x"80d0dc0c",
   693 => x"80d0f00c",
   694 => x"80d0e008",
   695 => x"80d0f408",
   696 => x"80d0e00c",
   697 => x"80d0f40c",
   698 => x"80d0e408",
   699 => x"80d0f808",
   700 => x"80d0e40c",
   701 => x"80d0f80c",
   702 => x"80d39408",
   703 => x"a0065280",
   704 => x"72259638",
   705 => x"91e52d8e",
   706 => x"832d80d0",
   707 => x"fc088132",
   708 => x"7080d0fc",
   709 => x"0c5185b2",
   710 => x"2d80d0fc",
   711 => x"0882ef38",
   712 => x"80d0e808",
   713 => x"518fca2d",
   714 => x"80d2bc08",
   715 => x"802e8b38",
   716 => x"80d39c08",
   717 => x"810780d3",
   718 => x"9c0c80d0",
   719 => x"ec08518f",
   720 => x"ca2d80d2",
   721 => x"bc08802e",
   722 => x"8b3880d3",
   723 => x"9c088207",
   724 => x"80d39c0c",
   725 => x"80d0f008",
   726 => x"518fca2d",
   727 => x"80d2bc08",
   728 => x"802e8b38",
   729 => x"80d39c08",
   730 => x"840780d3",
   731 => x"9c0c80d0",
   732 => x"f408518f",
   733 => x"ca2d80d2",
   734 => x"bc08802e",
   735 => x"8b3880d3",
   736 => x"9c088807",
   737 => x"80d39c0c",
   738 => x"80d0f808",
   739 => x"518fca2d",
   740 => x"80d2bc08",
   741 => x"802e8b38",
   742 => x"80d39c08",
   743 => x"900780d3",
   744 => x"9c0c80d0",
   745 => x"d408518f",
   746 => x"ca2d80d2",
   747 => x"bc08802e",
   748 => x"8c3880d3",
   749 => x"9c088280",
   750 => x"0780d39c",
   751 => x"0c80d0d8",
   752 => x"08518fca",
   753 => x"2d80d2bc",
   754 => x"08802e8c",
   755 => x"3880d39c",
   756 => x"08848007",
   757 => x"80d39c0c",
   758 => x"80d0dc08",
   759 => x"518fca2d",
   760 => x"80d2bc08",
   761 => x"802e8c38",
   762 => x"80d39c08",
   763 => x"88800780",
   764 => x"d39c0c80",
   765 => x"d0e00851",
   766 => x"8fca2d80",
   767 => x"d2bc0880",
   768 => x"2e8c3880",
   769 => x"d39c0890",
   770 => x"800780d3",
   771 => x"9c0c80d0",
   772 => x"e408518f",
   773 => x"ca2d80d2",
   774 => x"bc08802e",
   775 => x"8c3880d3",
   776 => x"9c08a080",
   777 => x"0780d39c",
   778 => x"0c94518f",
   779 => x"ca2d80d2",
   780 => x"bc085291",
   781 => x"518fca2d",
   782 => x"7180d2bc",
   783 => x"08065280",
   784 => x"e6518fca",
   785 => x"2d7180d2",
   786 => x"bc080652",
   787 => x"71802e8d",
   788 => x"3880d39c",
   789 => x"08848080",
   790 => x"0780d39c",
   791 => x"0c80fe51",
   792 => x"8fca2d80",
   793 => x"d2bc0852",
   794 => x"87518fca",
   795 => x"2d7180d2",
   796 => x"bc080752",
   797 => x"71802e8d",
   798 => x"3880d39c",
   799 => x"08888080",
   800 => x"0780d39c",
   801 => x"0c80d39c",
   802 => x"08ed0ca1",
   803 => x"99049451",
   804 => x"8fca2d80",
   805 => x"d2bc0852",
   806 => x"91518fca",
   807 => x"2d7180d2",
   808 => x"bc080652",
   809 => x"80e6518f",
   810 => x"ca2d7180",
   811 => x"d2bc0806",
   812 => x"5271802e",
   813 => x"8d3880d3",
   814 => x"9c088480",
   815 => x"800780d3",
   816 => x"9c0c80fe",
   817 => x"518fca2d",
   818 => x"80d2bc08",
   819 => x"5287518f",
   820 => x"ca2d7180",
   821 => x"d2bc0807",
   822 => x"5271802e",
   823 => x"8d3880d3",
   824 => x"9c088880",
   825 => x"800780d3",
   826 => x"9c0c80d3",
   827 => x"9c08ed0c",
   828 => x"81f5518f",
   829 => x"ca2d80d2",
   830 => x"bc08812a",
   831 => x"70810651",
   832 => x"5271a438",
   833 => x"80d0e808",
   834 => x"518fca2d",
   835 => x"80d2bc08",
   836 => x"812a7081",
   837 => x"06515271",
   838 => x"8e3880d3",
   839 => x"94088106",
   840 => x"52807225",
   841 => x"80c23880",
   842 => x"d3940881",
   843 => x"06528072",
   844 => x"25843891",
   845 => x"e52d80d3",
   846 => x"a8085271",
   847 => x"802e8a38",
   848 => x"ff1280d3",
   849 => x"a80c9ae8",
   850 => x"0480d3a4",
   851 => x"081080d3",
   852 => x"a4080570",
   853 => x"84291651",
   854 => x"52881208",
   855 => x"802e8938",
   856 => x"ff518812",
   857 => x"0852712d",
   858 => x"81f2518f",
   859 => x"ca2d80d2",
   860 => x"bc08812a",
   861 => x"70810651",
   862 => x"5271a438",
   863 => x"80d0ec08",
   864 => x"518fca2d",
   865 => x"80d2bc08",
   866 => x"812a7081",
   867 => x"06515271",
   868 => x"8e3880d3",
   869 => x"94088206",
   870 => x"52807225",
   871 => x"80c33880",
   872 => x"d3940882",
   873 => x"06528072",
   874 => x"25843891",
   875 => x"e52d80d3",
   876 => x"a408ff11",
   877 => x"80d3a808",
   878 => x"56535373",
   879 => x"72258a38",
   880 => x"811480d3",
   881 => x"a80c9be1",
   882 => x"04721013",
   883 => x"70842916",
   884 => x"51528812",
   885 => x"08802e89",
   886 => x"38fe5188",
   887 => x"12085271",
   888 => x"2d81fd51",
   889 => x"8fca2d80",
   890 => x"d2bc0881",
   891 => x"2a708106",
   892 => x"515271a4",
   893 => x"3880d0f0",
   894 => x"08518fca",
   895 => x"2d80d2bc",
   896 => x"08812a70",
   897 => x"81065152",
   898 => x"718e3880",
   899 => x"d3940884",
   900 => x"06528072",
   901 => x"2580c038",
   902 => x"80d39408",
   903 => x"84065280",
   904 => x"72258438",
   905 => x"91e52d80",
   906 => x"d3a80880",
   907 => x"2e8a3880",
   908 => x"0b80d3a8",
   909 => x"0c9cd704",
   910 => x"80d3a408",
   911 => x"1080d3a4",
   912 => x"08057084",
   913 => x"29165152",
   914 => x"88120880",
   915 => x"2e8938fd",
   916 => x"51881208",
   917 => x"52712d81",
   918 => x"fa518fca",
   919 => x"2d80d2bc",
   920 => x"08812a70",
   921 => x"81065152",
   922 => x"71a43880",
   923 => x"d0f40851",
   924 => x"8fca2d80",
   925 => x"d2bc0881",
   926 => x"2a708106",
   927 => x"5152718e",
   928 => x"3880d394",
   929 => x"08880652",
   930 => x"80722580",
   931 => x"c03880d3",
   932 => x"94088806",
   933 => x"52807225",
   934 => x"843891e5",
   935 => x"2d80d3a4",
   936 => x"08ff1154",
   937 => x"5280d3a8",
   938 => x"08732589",
   939 => x"387280d3",
   940 => x"a80c9dcd",
   941 => x"04711012",
   942 => x"70842916",
   943 => x"51528812",
   944 => x"08802e89",
   945 => x"38fc5188",
   946 => x"12085271",
   947 => x"2d80d3a8",
   948 => x"08705354",
   949 => x"73802e8a",
   950 => x"388c15ff",
   951 => x"1555559d",
   952 => x"d404820b",
   953 => x"80d2d00c",
   954 => x"718f0680",
   955 => x"d2cc0c81",
   956 => x"eb518fca",
   957 => x"2d80d2bc",
   958 => x"08812a70",
   959 => x"81065152",
   960 => x"71802ead",
   961 => x"38740885",
   962 => x"2e098106",
   963 => x"a4388815",
   964 => x"80f52dff",
   965 => x"05527188",
   966 => x"1681b72d",
   967 => x"71982b52",
   968 => x"71802588",
   969 => x"38800b88",
   970 => x"1681b72d",
   971 => x"745192de",
   972 => x"2d81f451",
   973 => x"8fca2d80",
   974 => x"d2bc0881",
   975 => x"2a708106",
   976 => x"51527180",
   977 => x"2eb33874",
   978 => x"08852e09",
   979 => x"8106aa38",
   980 => x"881580f5",
   981 => x"2d810552",
   982 => x"71881681",
   983 => x"b72d7181",
   984 => x"ff068b16",
   985 => x"80f52d54",
   986 => x"52727227",
   987 => x"87387288",
   988 => x"1681b72d",
   989 => x"745192de",
   990 => x"2d80da51",
   991 => x"8fca2d80",
   992 => x"d2bc0881",
   993 => x"2a708106",
   994 => x"5152718e",
   995 => x"3880d394",
   996 => x"08900652",
   997 => x"80722581",
   998 => x"bc3880d3",
   999 => x"a00880d3",
  1000 => x"94089006",
  1001 => x"53538072",
  1002 => x"25843891",
  1003 => x"e52d80d3",
  1004 => x"a8085473",
  1005 => x"802e8a38",
  1006 => x"8c13ff15",
  1007 => x"55539fb3",
  1008 => x"04720852",
  1009 => x"71822ea6",
  1010 => x"38718226",
  1011 => x"89387181",
  1012 => x"2eaa38a0",
  1013 => x"d5047183",
  1014 => x"2eb43871",
  1015 => x"842e0981",
  1016 => x"0680f238",
  1017 => x"88130851",
  1018 => x"94b42da0",
  1019 => x"d50480d3",
  1020 => x"a8085188",
  1021 => x"13085271",
  1022 => x"2da0d504",
  1023 => x"810b8814",
  1024 => x"082b80d0",
  1025 => x"d0083280",
  1026 => x"d0d00ca0",
  1027 => x"a9048813",
  1028 => x"80f52d81",
  1029 => x"058b1480",
  1030 => x"f52d5354",
  1031 => x"71742483",
  1032 => x"38805473",
  1033 => x"881481b7",
  1034 => x"2d938e2d",
  1035 => x"a0d50475",
  1036 => x"08802ea4",
  1037 => x"38750851",
  1038 => x"8fca2d80",
  1039 => x"d2bc0881",
  1040 => x"06527180",
  1041 => x"2e8c3880",
  1042 => x"d3a80851",
  1043 => x"84160852",
  1044 => x"712d8816",
  1045 => x"5675d838",
  1046 => x"8054800b",
  1047 => x"80d2d00c",
  1048 => x"738f0680",
  1049 => x"d2cc0ca0",
  1050 => x"527380d3",
  1051 => x"a8082e09",
  1052 => x"81069938",
  1053 => x"80d3a408",
  1054 => x"ff057432",
  1055 => x"70098105",
  1056 => x"7072079f",
  1057 => x"2a917131",
  1058 => x"51515353",
  1059 => x"71518384",
  1060 => x"2d811454",
  1061 => x"8e7425c2",
  1062 => x"3880d0fc",
  1063 => x"0880d2bc",
  1064 => x"0c029805",
  1065 => x"0d0402f4",
  1066 => x"050dd452",
  1067 => x"81ff720c",
  1068 => x"71085381",
  1069 => x"ff720c72",
  1070 => x"882b83fe",
  1071 => x"80067208",
  1072 => x"7081ff06",
  1073 => x"51525381",
  1074 => x"ff720c72",
  1075 => x"7107882b",
  1076 => x"72087081",
  1077 => x"ff065152",
  1078 => x"5381ff72",
  1079 => x"0c727107",
  1080 => x"882b7208",
  1081 => x"7081ff06",
  1082 => x"720780d2",
  1083 => x"bc0c5253",
  1084 => x"028c050d",
  1085 => x"0402f405",
  1086 => x"0d747671",
  1087 => x"81ff06d4",
  1088 => x"0c535380",
  1089 => x"d3b00885",
  1090 => x"3871892b",
  1091 => x"5271982a",
  1092 => x"d40c7190",
  1093 => x"2a7081ff",
  1094 => x"06d40c51",
  1095 => x"71882a70",
  1096 => x"81ff06d4",
  1097 => x"0c517181",
  1098 => x"ff06d40c",
  1099 => x"72902a70",
  1100 => x"81ff06d4",
  1101 => x"0c51d408",
  1102 => x"7081ff06",
  1103 => x"515182b8",
  1104 => x"bf527081",
  1105 => x"ff2e0981",
  1106 => x"06943881",
  1107 => x"ff0bd40c",
  1108 => x"d4087081",
  1109 => x"ff06ff14",
  1110 => x"54515171",
  1111 => x"e5387080",
  1112 => x"d2bc0c02",
  1113 => x"8c050d04",
  1114 => x"02fc050d",
  1115 => x"81c75181",
  1116 => x"ff0bd40c",
  1117 => x"ff115170",
  1118 => x"8025f438",
  1119 => x"0284050d",
  1120 => x"0402f405",
  1121 => x"0d81ff0b",
  1122 => x"d40c9353",
  1123 => x"805287fc",
  1124 => x"80c151a1",
  1125 => x"f52d80d2",
  1126 => x"bc088b38",
  1127 => x"81ff0bd4",
  1128 => x"0c8153a3",
  1129 => x"af04a2e8",
  1130 => x"2dff1353",
  1131 => x"72de3872",
  1132 => x"80d2bc0c",
  1133 => x"028c050d",
  1134 => x"0402ec05",
  1135 => x"0d810b80",
  1136 => x"d3b00c84",
  1137 => x"54d00870",
  1138 => x"8f2a7081",
  1139 => x"06515153",
  1140 => x"72f33872",
  1141 => x"d00ca2e8",
  1142 => x"2d80c8b4",
  1143 => x"5184a82d",
  1144 => x"d008708f",
  1145 => x"2a708106",
  1146 => x"51515372",
  1147 => x"f338810b",
  1148 => x"d00cb153",
  1149 => x"805284d4",
  1150 => x"80c051a1",
  1151 => x"f52d80d2",
  1152 => x"bc08812e",
  1153 => x"93387282",
  1154 => x"2ebf38ff",
  1155 => x"135372e4",
  1156 => x"38ff1454",
  1157 => x"73ffae38",
  1158 => x"a2e82d83",
  1159 => x"aa52849c",
  1160 => x"80c851a1",
  1161 => x"f52d80d2",
  1162 => x"bc08812e",
  1163 => x"09810693",
  1164 => x"38a1a62d",
  1165 => x"80d2bc08",
  1166 => x"83ffff06",
  1167 => x"537283aa",
  1168 => x"2e9f38a3",
  1169 => x"812da4dc",
  1170 => x"0480c8c0",
  1171 => x"5184a82d",
  1172 => x"8053a6b1",
  1173 => x"0480c8d8",
  1174 => x"5184a82d",
  1175 => x"8054a682",
  1176 => x"0481ff0b",
  1177 => x"d40cb154",
  1178 => x"a2e82d8f",
  1179 => x"cf538052",
  1180 => x"87fc80f7",
  1181 => x"51a1f52d",
  1182 => x"80d2bc08",
  1183 => x"5580d2bc",
  1184 => x"08812e09",
  1185 => x"81069c38",
  1186 => x"81ff0bd4",
  1187 => x"0c820a52",
  1188 => x"849c80e9",
  1189 => x"51a1f52d",
  1190 => x"80d2bc08",
  1191 => x"802e8d38",
  1192 => x"a2e82dff",
  1193 => x"135372c6",
  1194 => x"38a5f504",
  1195 => x"81ff0bd4",
  1196 => x"0c80d2bc",
  1197 => x"085287fc",
  1198 => x"80fa51a1",
  1199 => x"f52d80d2",
  1200 => x"bc08b238",
  1201 => x"81ff0bd4",
  1202 => x"0cd40853",
  1203 => x"81ff0bd4",
  1204 => x"0c81ff0b",
  1205 => x"d40c81ff",
  1206 => x"0bd40c81",
  1207 => x"ff0bd40c",
  1208 => x"72862a70",
  1209 => x"81067656",
  1210 => x"51537296",
  1211 => x"3880d2bc",
  1212 => x"0854a682",
  1213 => x"0473822e",
  1214 => x"fedb38ff",
  1215 => x"145473fe",
  1216 => x"e7387380",
  1217 => x"d3b00c73",
  1218 => x"8b388152",
  1219 => x"87fc80d0",
  1220 => x"51a1f52d",
  1221 => x"81ff0bd4",
  1222 => x"0cd00870",
  1223 => x"8f2a7081",
  1224 => x"06515153",
  1225 => x"72f33872",
  1226 => x"d00c81ff",
  1227 => x"0bd40c81",
  1228 => x"537280d2",
  1229 => x"bc0c0294",
  1230 => x"050d0402",
  1231 => x"e8050d78",
  1232 => x"55805681",
  1233 => x"ff0bd40c",
  1234 => x"d008708f",
  1235 => x"2a708106",
  1236 => x"51515372",
  1237 => x"f3388281",
  1238 => x"0bd00c81",
  1239 => x"ff0bd40c",
  1240 => x"775287fc",
  1241 => x"80d151a1",
  1242 => x"f52d80db",
  1243 => x"c6df5480",
  1244 => x"d2bc0880",
  1245 => x"2e8b3880",
  1246 => x"c8f85184",
  1247 => x"a82da7d5",
  1248 => x"0481ff0b",
  1249 => x"d40cd408",
  1250 => x"7081ff06",
  1251 => x"51537281",
  1252 => x"fe2e0981",
  1253 => x"069e3880",
  1254 => x"ff53a1a6",
  1255 => x"2d80d2bc",
  1256 => x"08757084",
  1257 => x"05570cff",
  1258 => x"13537280",
  1259 => x"25ec3881",
  1260 => x"56a7ba04",
  1261 => x"ff145473",
  1262 => x"c83881ff",
  1263 => x"0bd40c81",
  1264 => x"ff0bd40c",
  1265 => x"d008708f",
  1266 => x"2a708106",
  1267 => x"51515372",
  1268 => x"f33872d0",
  1269 => x"0c7580d2",
  1270 => x"bc0c0298",
  1271 => x"050d0402",
  1272 => x"e8050d77",
  1273 => x"797b5855",
  1274 => x"55805372",
  1275 => x"7625a338",
  1276 => x"74708105",
  1277 => x"5680f52d",
  1278 => x"74708105",
  1279 => x"5680f52d",
  1280 => x"52527171",
  1281 => x"2e863881",
  1282 => x"51a89404",
  1283 => x"811353a7",
  1284 => x"eb048051",
  1285 => x"7080d2bc",
  1286 => x"0c029805",
  1287 => x"0d0402ec",
  1288 => x"050d7655",
  1289 => x"74802e80",
  1290 => x"c2389a15",
  1291 => x"80e02d51",
  1292 => x"b6d92d80",
  1293 => x"d2bc0880",
  1294 => x"d2bc0880",
  1295 => x"d9e40c80",
  1296 => x"d2bc0854",
  1297 => x"5480d9c0",
  1298 => x"08802e9a",
  1299 => x"38941580",
  1300 => x"e02d51b6",
  1301 => x"d92d80d2",
  1302 => x"bc08902b",
  1303 => x"83fff00a",
  1304 => x"06707507",
  1305 => x"51537280",
  1306 => x"d9e40c80",
  1307 => x"d9e40853",
  1308 => x"72802e9d",
  1309 => x"3880d9b8",
  1310 => x"08fe1471",
  1311 => x"2980d9cc",
  1312 => x"080580d9",
  1313 => x"e80c7084",
  1314 => x"2b80d9c4",
  1315 => x"0c54a9bf",
  1316 => x"0480d9d0",
  1317 => x"0880d9e4",
  1318 => x"0c80d9d4",
  1319 => x"0880d9e8",
  1320 => x"0c80d9c0",
  1321 => x"08802e8b",
  1322 => x"3880d9b8",
  1323 => x"08842b53",
  1324 => x"a9ba0480",
  1325 => x"d9d80884",
  1326 => x"2b537280",
  1327 => x"d9c40c02",
  1328 => x"94050d04",
  1329 => x"02d8050d",
  1330 => x"800b80d9",
  1331 => x"c00c8454",
  1332 => x"a3b92d80",
  1333 => x"d2bc0880",
  1334 => x"2e973880",
  1335 => x"d3b45280",
  1336 => x"51a6bb2d",
  1337 => x"80d2bc08",
  1338 => x"802e8638",
  1339 => x"fe54a9f9",
  1340 => x"04ff1454",
  1341 => x"738024d8",
  1342 => x"38738d38",
  1343 => x"80c98851",
  1344 => x"84a82d73",
  1345 => x"55afce04",
  1346 => x"8056810b",
  1347 => x"80d9ec0c",
  1348 => x"885380c9",
  1349 => x"9c5280d3",
  1350 => x"ea51a7df",
  1351 => x"2d80d2bc",
  1352 => x"08762e09",
  1353 => x"81068938",
  1354 => x"80d2bc08",
  1355 => x"80d9ec0c",
  1356 => x"885380c9",
  1357 => x"a85280d4",
  1358 => x"8651a7df",
  1359 => x"2d80d2bc",
  1360 => x"08893880",
  1361 => x"d2bc0880",
  1362 => x"d9ec0c80",
  1363 => x"d9ec0880",
  1364 => x"2e818138",
  1365 => x"80d6fa0b",
  1366 => x"80f52d80",
  1367 => x"d6fb0b80",
  1368 => x"f52d7198",
  1369 => x"2b71902b",
  1370 => x"0780d6fc",
  1371 => x"0b80f52d",
  1372 => x"70882b72",
  1373 => x"0780d6fd",
  1374 => x"0b80f52d",
  1375 => x"710780d7",
  1376 => x"b20b80f5",
  1377 => x"2d80d7b3",
  1378 => x"0b80f52d",
  1379 => x"71882b07",
  1380 => x"535f5452",
  1381 => x"5a565755",
  1382 => x"7381abaa",
  1383 => x"2e098106",
  1384 => x"8e387551",
  1385 => x"b6a82d80",
  1386 => x"d2bc0856",
  1387 => x"abbd0473",
  1388 => x"82d4d52e",
  1389 => x"883880c9",
  1390 => x"b451ac89",
  1391 => x"0480d3b4",
  1392 => x"527551a6",
  1393 => x"bb2d80d2",
  1394 => x"bc085580",
  1395 => x"d2bc0880",
  1396 => x"2e83fb38",
  1397 => x"885380c9",
  1398 => x"a85280d4",
  1399 => x"8651a7df",
  1400 => x"2d80d2bc",
  1401 => x"088a3881",
  1402 => x"0b80d9c0",
  1403 => x"0cac8f04",
  1404 => x"885380c9",
  1405 => x"9c5280d3",
  1406 => x"ea51a7df",
  1407 => x"2d80d2bc",
  1408 => x"08802e8b",
  1409 => x"3880c9c8",
  1410 => x"5184a82d",
  1411 => x"acee0480",
  1412 => x"d7b20b80",
  1413 => x"f52d5473",
  1414 => x"80d52e09",
  1415 => x"810680ce",
  1416 => x"3880d7b3",
  1417 => x"0b80f52d",
  1418 => x"547381aa",
  1419 => x"2e098106",
  1420 => x"bd38800b",
  1421 => x"80d3b40b",
  1422 => x"80f52d56",
  1423 => x"547481e9",
  1424 => x"2e833881",
  1425 => x"547481eb",
  1426 => x"2e8c3880",
  1427 => x"5573752e",
  1428 => x"09810682",
  1429 => x"f93880d3",
  1430 => x"bf0b80f5",
  1431 => x"2d55748e",
  1432 => x"3880d3c0",
  1433 => x"0b80f52d",
  1434 => x"5473822e",
  1435 => x"86388055",
  1436 => x"afce0480",
  1437 => x"d3c10b80",
  1438 => x"f52d7080",
  1439 => x"d9b80cff",
  1440 => x"0580d9bc",
  1441 => x"0c80d3c2",
  1442 => x"0b80f52d",
  1443 => x"80d3c30b",
  1444 => x"80f52d58",
  1445 => x"76057782",
  1446 => x"80290570",
  1447 => x"80d9c80c",
  1448 => x"80d3c40b",
  1449 => x"80f52d70",
  1450 => x"80d9dc0c",
  1451 => x"80d9c008",
  1452 => x"59575876",
  1453 => x"802e81b7",
  1454 => x"38885380",
  1455 => x"c9a85280",
  1456 => x"d48651a7",
  1457 => x"df2d80d2",
  1458 => x"bc088282",
  1459 => x"3880d9b8",
  1460 => x"0870842b",
  1461 => x"80d9c40c",
  1462 => x"7080d9d8",
  1463 => x"0c80d3d9",
  1464 => x"0b80f52d",
  1465 => x"80d3d80b",
  1466 => x"80f52d71",
  1467 => x"82802905",
  1468 => x"80d3da0b",
  1469 => x"80f52d70",
  1470 => x"84808029",
  1471 => x"1280d3db",
  1472 => x"0b80f52d",
  1473 => x"7081800a",
  1474 => x"29127080",
  1475 => x"d9e00c80",
  1476 => x"d9dc0871",
  1477 => x"2980d9c8",
  1478 => x"08057080",
  1479 => x"d9cc0c80",
  1480 => x"d3e10b80",
  1481 => x"f52d80d3",
  1482 => x"e00b80f5",
  1483 => x"2d718280",
  1484 => x"290580d3",
  1485 => x"e20b80f5",
  1486 => x"2d708480",
  1487 => x"80291280",
  1488 => x"d3e30b80",
  1489 => x"f52d7098",
  1490 => x"2b81f00a",
  1491 => x"06720570",
  1492 => x"80d9d00c",
  1493 => x"fe117e29",
  1494 => x"770580d9",
  1495 => x"d40c5259",
  1496 => x"5243545e",
  1497 => x"51525952",
  1498 => x"5d575957",
  1499 => x"afc70480",
  1500 => x"d3c60b80",
  1501 => x"f52d80d3",
  1502 => x"c50b80f5",
  1503 => x"2d718280",
  1504 => x"29057080",
  1505 => x"d9c40c70",
  1506 => x"a02983ff",
  1507 => x"0570892a",
  1508 => x"7080d9d8",
  1509 => x"0c80d3cb",
  1510 => x"0b80f52d",
  1511 => x"80d3ca0b",
  1512 => x"80f52d71",
  1513 => x"82802905",
  1514 => x"7080d9e0",
  1515 => x"0c7b7129",
  1516 => x"1e7080d9",
  1517 => x"d40c7d80",
  1518 => x"d9d00c73",
  1519 => x"0580d9cc",
  1520 => x"0c555e51",
  1521 => x"51555580",
  1522 => x"51a89e2d",
  1523 => x"81557480",
  1524 => x"d2bc0c02",
  1525 => x"a8050d04",
  1526 => x"02ec050d",
  1527 => x"7670872c",
  1528 => x"7180ff06",
  1529 => x"55565480",
  1530 => x"d9c0088a",
  1531 => x"3873882c",
  1532 => x"7481ff06",
  1533 => x"545580d3",
  1534 => x"b45280d9",
  1535 => x"c8081551",
  1536 => x"a6bb2d80",
  1537 => x"d2bc0854",
  1538 => x"80d2bc08",
  1539 => x"802eb838",
  1540 => x"80d9c008",
  1541 => x"802e9a38",
  1542 => x"72842980",
  1543 => x"d3b40570",
  1544 => x"085253b6",
  1545 => x"a82d80d2",
  1546 => x"bc08f00a",
  1547 => x"0653b0c5",
  1548 => x"04721080",
  1549 => x"d3b40570",
  1550 => x"80e02d52",
  1551 => x"53b6d92d",
  1552 => x"80d2bc08",
  1553 => x"53725473",
  1554 => x"80d2bc0c",
  1555 => x"0294050d",
  1556 => x"0402e005",
  1557 => x"0d797084",
  1558 => x"2c80d9e8",
  1559 => x"0805718f",
  1560 => x"06525553",
  1561 => x"728a3880",
  1562 => x"d3b45273",
  1563 => x"51a6bb2d",
  1564 => x"72a02980",
  1565 => x"d3b40554",
  1566 => x"807480f5",
  1567 => x"2d565374",
  1568 => x"732e8338",
  1569 => x"81537481",
  1570 => x"e52e81f4",
  1571 => x"38817074",
  1572 => x"06545872",
  1573 => x"802e81e8",
  1574 => x"388b1480",
  1575 => x"f52d7083",
  1576 => x"2a790658",
  1577 => x"56769b38",
  1578 => x"80d18008",
  1579 => x"53728938",
  1580 => x"7280d7b4",
  1581 => x"0b81b72d",
  1582 => x"7680d180",
  1583 => x"0c7353b3",
  1584 => x"8204758f",
  1585 => x"2e098106",
  1586 => x"81b63874",
  1587 => x"9f068d29",
  1588 => x"80d7a711",
  1589 => x"51538114",
  1590 => x"80f52d73",
  1591 => x"70810555",
  1592 => x"81b72d83",
  1593 => x"1480f52d",
  1594 => x"73708105",
  1595 => x"5581b72d",
  1596 => x"851480f5",
  1597 => x"2d737081",
  1598 => x"055581b7",
  1599 => x"2d871480",
  1600 => x"f52d7370",
  1601 => x"81055581",
  1602 => x"b72d8914",
  1603 => x"80f52d73",
  1604 => x"70810555",
  1605 => x"81b72d8e",
  1606 => x"1480f52d",
  1607 => x"73708105",
  1608 => x"5581b72d",
  1609 => x"901480f5",
  1610 => x"2d737081",
  1611 => x"055581b7",
  1612 => x"2d921480",
  1613 => x"f52d7370",
  1614 => x"81055581",
  1615 => x"b72d9414",
  1616 => x"80f52d73",
  1617 => x"70810555",
  1618 => x"81b72d96",
  1619 => x"1480f52d",
  1620 => x"73708105",
  1621 => x"5581b72d",
  1622 => x"981480f5",
  1623 => x"2d737081",
  1624 => x"055581b7",
  1625 => x"2d9c1480",
  1626 => x"f52d7370",
  1627 => x"81055581",
  1628 => x"b72d9e14",
  1629 => x"80f52d73",
  1630 => x"81b72d77",
  1631 => x"80d1800c",
  1632 => x"80537280",
  1633 => x"d2bc0c02",
  1634 => x"a0050d04",
  1635 => x"02cc050d",
  1636 => x"7e605e5b",
  1637 => x"800b80d9",
  1638 => x"e40880d9",
  1639 => x"e808595d",
  1640 => x"56805980",
  1641 => x"d9c40879",
  1642 => x"2e81de38",
  1643 => x"788f06a0",
  1644 => x"17575473",
  1645 => x"913880d3",
  1646 => x"b4527651",
  1647 => x"811757a6",
  1648 => x"bb2d80d3",
  1649 => x"b4568076",
  1650 => x"80f52d56",
  1651 => x"5474742e",
  1652 => x"83388154",
  1653 => x"7481e52e",
  1654 => x"81a33881",
  1655 => x"70750655",
  1656 => x"5a73802e",
  1657 => x"8197388b",
  1658 => x"1680f52d",
  1659 => x"70980659",
  1660 => x"547780e3",
  1661 => x"388b537c",
  1662 => x"527551a7",
  1663 => x"df2d80d2",
  1664 => x"bc0880f9",
  1665 => x"389c1608",
  1666 => x"51b6a82d",
  1667 => x"80d2bc08",
  1668 => x"841c0c9a",
  1669 => x"1680e02d",
  1670 => x"51b6d92d",
  1671 => x"80d2bc08",
  1672 => x"80d2bc08",
  1673 => x"881d0c80",
  1674 => x"d2bc0855",
  1675 => x"5580d9c0",
  1676 => x"08802e99",
  1677 => x"38941680",
  1678 => x"e02d51b6",
  1679 => x"d92d80d2",
  1680 => x"bc08902b",
  1681 => x"83fff00a",
  1682 => x"06701651",
  1683 => x"5473881c",
  1684 => x"0c777b0c",
  1685 => x"b4f80473",
  1686 => x"842a7081",
  1687 => x"06515473",
  1688 => x"802e9a38",
  1689 => x"8b537c52",
  1690 => x"7551a7df",
  1691 => x"2d80d2bc",
  1692 => x"088b3875",
  1693 => x"51a89e2d",
  1694 => x"7954b5c5",
  1695 => x"04811959",
  1696 => x"80d9c408",
  1697 => x"7926fea4",
  1698 => x"3880d9c0",
  1699 => x"08802eb3",
  1700 => x"387b51af",
  1701 => x"d82d80d2",
  1702 => x"bc0880d2",
  1703 => x"bc0880ff",
  1704 => x"fffff806",
  1705 => x"555c7380",
  1706 => x"fffffff8",
  1707 => x"2e953880",
  1708 => x"d2bc08fe",
  1709 => x"0580d9b8",
  1710 => x"082980d9",
  1711 => x"cc080557",
  1712 => x"b3a10480",
  1713 => x"547380d2",
  1714 => x"bc0c02b4",
  1715 => x"050d0402",
  1716 => x"f4050d74",
  1717 => x"70088105",
  1718 => x"710c7008",
  1719 => x"80d9bc08",
  1720 => x"06535371",
  1721 => x"8f388813",
  1722 => x"0851afd8",
  1723 => x"2d80d2bc",
  1724 => x"0888140c",
  1725 => x"810b80d2",
  1726 => x"bc0c028c",
  1727 => x"050d0402",
  1728 => x"f0050d75",
  1729 => x"881108fe",
  1730 => x"0580d9b8",
  1731 => x"082980d9",
  1732 => x"cc081172",
  1733 => x"0880d9bc",
  1734 => x"08060579",
  1735 => x"55535454",
  1736 => x"a6bb2d02",
  1737 => x"90050d04",
  1738 => x"02f4050d",
  1739 => x"7470882a",
  1740 => x"83fe8006",
  1741 => x"7072982a",
  1742 => x"0772882b",
  1743 => x"87fc8080",
  1744 => x"0673982b",
  1745 => x"81f00a06",
  1746 => x"71730707",
  1747 => x"80d2bc0c",
  1748 => x"56515351",
  1749 => x"028c050d",
  1750 => x"0402f805",
  1751 => x"0d028e05",
  1752 => x"80f52d74",
  1753 => x"882b0770",
  1754 => x"83ffff06",
  1755 => x"80d2bc0c",
  1756 => x"51028805",
  1757 => x"0d0402f4",
  1758 => x"050d7476",
  1759 => x"78535452",
  1760 => x"80712597",
  1761 => x"38727081",
  1762 => x"055480f5",
  1763 => x"2d727081",
  1764 => x"055481b7",
  1765 => x"2dff1151",
  1766 => x"70eb3880",
  1767 => x"7281b72d",
  1768 => x"028c050d",
  1769 => x"0402e805",
  1770 => x"0d775680",
  1771 => x"70565473",
  1772 => x"7624b638",
  1773 => x"80d9c408",
  1774 => x"742eae38",
  1775 => x"7351b0d1",
  1776 => x"2d80d2bc",
  1777 => x"0880d2bc",
  1778 => x"08098105",
  1779 => x"7080d2bc",
  1780 => x"08079f2a",
  1781 => x"77058117",
  1782 => x"57575353",
  1783 => x"74762489",
  1784 => x"3880d9c4",
  1785 => x"087426d4",
  1786 => x"387280d2",
  1787 => x"bc0c0298",
  1788 => x"050d0402",
  1789 => x"f0050d80",
  1790 => x"d2b80816",
  1791 => x"51b7a52d",
  1792 => x"80d2bc08",
  1793 => x"802e9f38",
  1794 => x"8b5380d2",
  1795 => x"bc085280",
  1796 => x"d7b451b6",
  1797 => x"f62d80d9",
  1798 => x"f0085473",
  1799 => x"802e8738",
  1800 => x"80d7b451",
  1801 => x"732d0290",
  1802 => x"050d0402",
  1803 => x"dc050d80",
  1804 => x"705a5574",
  1805 => x"80d2b808",
  1806 => x"25b43880",
  1807 => x"d9c40875",
  1808 => x"2eac3878",
  1809 => x"51b0d12d",
  1810 => x"80d2bc08",
  1811 => x"09810570",
  1812 => x"80d2bc08",
  1813 => x"079f2a76",
  1814 => x"05811b5b",
  1815 => x"56547480",
  1816 => x"d2b80825",
  1817 => x"893880d9",
  1818 => x"c4087926",
  1819 => x"d6388055",
  1820 => x"7880d9c4",
  1821 => x"082781db",
  1822 => x"387851b0",
  1823 => x"d12d80d2",
  1824 => x"bc08802e",
  1825 => x"81ad3880",
  1826 => x"d2bc088b",
  1827 => x"0580f52d",
  1828 => x"70842a70",
  1829 => x"81067710",
  1830 => x"78842b80",
  1831 => x"d7b40b80",
  1832 => x"f52d5c5c",
  1833 => x"53515556",
  1834 => x"73802e80",
  1835 => x"cb387416",
  1836 => x"822bbaf7",
  1837 => x"0b80d18c",
  1838 => x"120c5477",
  1839 => x"75311080",
  1840 => x"d9f41155",
  1841 => x"56907470",
  1842 => x"81055681",
  1843 => x"b72da074",
  1844 => x"81b72d76",
  1845 => x"81ff0681",
  1846 => x"16585473",
  1847 => x"802e8a38",
  1848 => x"9c5380d7",
  1849 => x"b452b9f0",
  1850 => x"048b5380",
  1851 => x"d2bc0852",
  1852 => x"80d9f616",
  1853 => x"51baab04",
  1854 => x"7416822b",
  1855 => x"b7f30b80",
  1856 => x"d18c120c",
  1857 => x"547681ff",
  1858 => x"06811658",
  1859 => x"5473802e",
  1860 => x"8a389c53",
  1861 => x"80d7b452",
  1862 => x"baa2048b",
  1863 => x"5380d2bc",
  1864 => x"08527775",
  1865 => x"311080d9",
  1866 => x"f4055176",
  1867 => x"55b6f62d",
  1868 => x"bac80474",
  1869 => x"90297531",
  1870 => x"701080d9",
  1871 => x"f4055154",
  1872 => x"80d2bc08",
  1873 => x"7481b72d",
  1874 => x"81195974",
  1875 => x"8b24a338",
  1876 => x"b8f00474",
  1877 => x"90297531",
  1878 => x"701080d9",
  1879 => x"f4058c77",
  1880 => x"31575154",
  1881 => x"807481b7",
  1882 => x"2d9e14ff",
  1883 => x"16565474",
  1884 => x"f33802a4",
  1885 => x"050d0402",
  1886 => x"fc050d80",
  1887 => x"d2b80813",
  1888 => x"51b7a52d",
  1889 => x"80d2bc08",
  1890 => x"802e8938",
  1891 => x"80d2bc08",
  1892 => x"51a89e2d",
  1893 => x"800b80d2",
  1894 => x"b80cb8ab",
  1895 => x"2d938e2d",
  1896 => x"0284050d",
  1897 => x"0402fc05",
  1898 => x"0d725170",
  1899 => x"fd2eb038",
  1900 => x"70fd248a",
  1901 => x"3870fc2e",
  1902 => x"80cc38bc",
  1903 => x"900470fe",
  1904 => x"2eb73870",
  1905 => x"ff2e0981",
  1906 => x"0680c538",
  1907 => x"80d2b808",
  1908 => x"5170802e",
  1909 => x"bb38ff11",
  1910 => x"80d2b80c",
  1911 => x"bc900480",
  1912 => x"d2b808f4",
  1913 => x"057080d2",
  1914 => x"b80c5170",
  1915 => x"8025a138",
  1916 => x"800b80d2",
  1917 => x"b80cbc90",
  1918 => x"0480d2b8",
  1919 => x"08810580",
  1920 => x"d2b80cbc",
  1921 => x"900480d2",
  1922 => x"b8088c05",
  1923 => x"80d2b80c",
  1924 => x"b8ab2d93",
  1925 => x"8e2d0284",
  1926 => x"050d0402",
  1927 => x"fc050d80",
  1928 => x"0b80d2b8",
  1929 => x"0cb8ab2d",
  1930 => x"91fc2d80",
  1931 => x"d2bc0880",
  1932 => x"d2a80c80",
  1933 => x"d1845194",
  1934 => x"b42d0284",
  1935 => x"050d0402",
  1936 => x"f8050d80",
  1937 => x"d2e408bf",
  1938 => x"f9ff0681",
  1939 => x"80077080",
  1940 => x"d2e40cfc",
  1941 => x"0c7351bc",
  1942 => x"9b2d0288",
  1943 => x"050d0402",
  1944 => x"f8050d80",
  1945 => x"d2e408bf",
  1946 => x"ffff0687",
  1947 => x"80077080",
  1948 => x"d2e40cfc",
  1949 => x"0c7351bc",
  1950 => x"9b2d0288",
  1951 => x"050d0471",
  1952 => x"80d9f00c",
  1953 => x"04000000",
  1954 => x"00ffffff",
  1955 => x"ff00ffff",
  1956 => x"ffff00ff",
  1957 => x"ffffff00",
  1958 => x"436f6e74",
  1959 => x"696e7565",
  1960 => x"00000000",
  1961 => x"3d205a58",
  1962 => x"38312f5a",
  1963 => x"58383020",
  1964 => x"436f6e66",
  1965 => x"69677572",
  1966 => x"6174696f",
  1967 => x"6e203d00",
  1968 => x"3d3d3d3d",
  1969 => x"3d3d3d3d",
  1970 => x"3d3d3d3d",
  1971 => x"3d3d3d3d",
  1972 => x"3d3d3d3d",
  1973 => x"3d3d3d3d",
  1974 => x"3d3d3d00",
  1975 => x"4c6f7720",
  1976 => x"52414d3a",
  1977 => x"204f6666",
  1978 => x"2f384b42",
  1979 => x"00000000",
  1980 => x"51532043",
  1981 => x"4852533a",
  1982 => x"44697361",
  1983 => x"626c6564",
  1984 => x"2f456e61",
  1985 => x"626c6564",
  1986 => x"28463129",
  1987 => x"00000000",
  1988 => x"4348524f",
  1989 => x"4d413831",
  1990 => x"3a204469",
  1991 => x"7361626c",
  1992 => x"65642f45",
  1993 => x"6e61626c",
  1994 => x"65640000",
  1995 => x"496e7665",
  1996 => x"72736520",
  1997 => x"76696465",
  1998 => x"6f3a204f",
  1999 => x"66662f4f",
  2000 => x"6e000000",
  2001 => x"426c6163",
  2002 => x"6b20626f",
  2003 => x"72646572",
  2004 => x"3a204f66",
  2005 => x"662f4f6e",
  2006 => x"00000000",
  2007 => x"56696465",
  2008 => x"6f206672",
  2009 => x"65717565",
  2010 => x"6e63793a",
  2011 => x"20353048",
  2012 => x"7a2f3630",
  2013 => x"487a0000",
  2014 => x"476f2042",
  2015 => x"61636b00",
  2016 => x"536c6f77",
  2017 => x"206d6f64",
  2018 => x"65207370",
  2019 => x"6565643a",
  2020 => x"204f7269",
  2021 => x"67696e61",
  2022 => x"6c000000",
  2023 => x"536c6f77",
  2024 => x"206d6f64",
  2025 => x"65207370",
  2026 => x"6565643a",
  2027 => x"204e6f57",
  2028 => x"61697400",
  2029 => x"536c6f77",
  2030 => x"206d6f64",
  2031 => x"65207370",
  2032 => x"6565643a",
  2033 => x"20783200",
  2034 => x"536c6f77",
  2035 => x"206d6f64",
  2036 => x"65207370",
  2037 => x"6565643a",
  2038 => x"20783800",
  2039 => x"43485224",
  2040 => x"3132382f",
  2041 => x"5544473a",
  2042 => x"20313238",
  2043 => x"20436861",
  2044 => x"72730000",
  2045 => x"43485224",
  2046 => x"3132382f",
  2047 => x"5544473a",
  2048 => x"20363420",
  2049 => x"43686172",
  2050 => x"73000000",
  2051 => x"43485224",
  2052 => x"3132382f",
  2053 => x"5544473a",
  2054 => x"20446973",
  2055 => x"61626c65",
  2056 => x"64000000",
  2057 => x"4a6f7973",
  2058 => x"7469636b",
  2059 => x"3a204375",
  2060 => x"72736f72",
  2061 => x"00000000",
  2062 => x"4a6f7973",
  2063 => x"7469636b",
  2064 => x"3a205369",
  2065 => x"6e636c61",
  2066 => x"69720000",
  2067 => x"4a6f7973",
  2068 => x"7469636b",
  2069 => x"3a205a58",
  2070 => x"38310000",
  2071 => x"4d61696e",
  2072 => x"2052414d",
  2073 => x"3a203136",
  2074 => x"4b420000",
  2075 => x"4d61696e",
  2076 => x"2052414d",
  2077 => x"3a203332",
  2078 => x"4b420000",
  2079 => x"4d61696e",
  2080 => x"2052414d",
  2081 => x"3a203438",
  2082 => x"4b420000",
  2083 => x"4d61696e",
  2084 => x"2052414d",
  2085 => x"3a20314b",
  2086 => x"42000000",
  2087 => x"436f6d70",
  2088 => x"75746572",
  2089 => x"204d6f64",
  2090 => x"656c3a20",
  2091 => x"5a583831",
  2092 => x"00000000",
  2093 => x"436f6d70",
  2094 => x"75746572",
  2095 => x"204d6f64",
  2096 => x"656c3a20",
  2097 => x"5a583830",
  2098 => x"00000000",
  2099 => x"3d3d205a",
  2100 => x"5838312f",
  2101 => x"5a583830",
  2102 => x"20666f72",
  2103 => x"205a5844",
  2104 => x"4f53203d",
  2105 => x"3d000000",
  2106 => x"3d3d3d3d",
  2107 => x"3d3d3d3d",
  2108 => x"3d3d3d3d",
  2109 => x"3d3d3d3d",
  2110 => x"3d3d3d3d",
  2111 => x"3d3d3d3d",
  2112 => x"3d000000",
  2113 => x"52657365",
  2114 => x"74000000",
  2115 => x"4c6f6164",
  2116 => x"20546170",
  2117 => x"6520282e",
  2118 => x"70292010",
  2119 => x"00000000",
  2120 => x"4c6f6164",
  2121 => x"20526f6d",
  2122 => x"2020282e",
  2123 => x"726f6d29",
  2124 => x"20100000",
  2125 => x"436f6e66",
  2126 => x"69677572",
  2127 => x"6174696f",
  2128 => x"6e206f70",
  2129 => x"74696f6e",
  2130 => x"73201000",
  2131 => x"4b657962",
  2132 => x"6f617264",
  2133 => x"2048656c",
  2134 => x"70000000",
  2135 => x"45786974",
  2136 => x"00000000",
  2137 => x"524f4d20",
  2138 => x"6c6f6164",
  2139 => x"696e6720",
  2140 => x"6661696c",
  2141 => x"65640000",
  2142 => x"4f4b0000",
  2143 => x"54617065",
  2144 => x"2066696c",
  2145 => x"65204c6f",
  2146 => x"61646564",
  2147 => x"2e000000",
  2148 => x"54797065",
  2149 => x"204c4f41",
  2150 => x"44202222",
  2151 => x"202b2045",
  2152 => x"4e544552",
  2153 => x"206f6e20",
  2154 => x"5a583831",
  2155 => x"00000000",
  2156 => x"5468656e",
  2157 => x"20707265",
  2158 => x"73732050",
  2159 => x"6c617920",
  2160 => x"616e6420",
  2161 => x"77616974",
  2162 => x"00000000",
  2163 => x"54686572",
  2164 => x"65206973",
  2165 => x"206e6f20",
  2166 => x"696d6167",
  2167 => x"65207768",
  2168 => x"656e206c",
  2169 => x"6f616469",
  2170 => x"6e670000",
  2171 => x"4c6f6164",
  2172 => x"20546170",
  2173 => x"6520282e",
  2174 => x"702c202e",
  2175 => x"38312920",
  2176 => x"10000000",
  2177 => x"3d205a58",
  2178 => x"38312f5a",
  2179 => x"58383020",
  2180 => x"4b657962",
  2181 => x"6f617264",
  2182 => x"2048656c",
  2183 => x"70203d00",
  2184 => x"5363726f",
  2185 => x"6c6c204c",
  2186 => x"6f636b3a",
  2187 => x"20636861",
  2188 => x"6e676520",
  2189 => x"62657477",
  2190 => x"65656e00",
  2191 => x"52474220",
  2192 => x"616e6420",
  2193 => x"56474120",
  2194 => x"76696465",
  2195 => x"6f206d6f",
  2196 => x"64650000",
  2197 => x"4374726c",
  2198 => x"2b416c74",
  2199 => x"2b44656c",
  2200 => x"6574653a",
  2201 => x"20536f66",
  2202 => x"74205265",
  2203 => x"73657400",
  2204 => x"4374726c",
  2205 => x"2b416c74",
  2206 => x"2b426163",
  2207 => x"6b737061",
  2208 => x"63653a20",
  2209 => x"48617264",
  2210 => x"20726573",
  2211 => x"65740000",
  2212 => x"45736320",
  2213 => x"6f72206a",
  2214 => x"6f797374",
  2215 => x"69636b20",
  2216 => x"62742e32",
  2217 => x"3a20746f",
  2218 => x"2073686f",
  2219 => x"77000000",
  2220 => x"6f722068",
  2221 => x"69646520",
  2222 => x"74686520",
  2223 => x"6f707469",
  2224 => x"6f6e7320",
  2225 => x"6d656e75",
  2226 => x"2e000000",
  2227 => x"57415344",
  2228 => x"202f2063",
  2229 => x"7572736f",
  2230 => x"72206b65",
  2231 => x"7973202f",
  2232 => x"206a6f79",
  2233 => x"73746963",
  2234 => x"6b000000",
  2235 => x"746f2073",
  2236 => x"656c6563",
  2237 => x"74206d65",
  2238 => x"6e75206f",
  2239 => x"7074696f",
  2240 => x"6e2e0000",
  2241 => x"456e7465",
  2242 => x"72202f20",
  2243 => x"46697265",
  2244 => x"20746f20",
  2245 => x"63686f6f",
  2246 => x"7365206f",
  2247 => x"7074696f",
  2248 => x"6e2e0000",
  2249 => x"3d205a58",
  2250 => x"38312f5a",
  2251 => x"58383020",
  2252 => x"436f7265",
  2253 => x"20437265",
  2254 => x"64697473",
  2255 => x"20203d00",
  2256 => x"43686970",
  2257 => x"2d382063",
  2258 => x"6f726520",
  2259 => x"666f7220",
  2260 => x"5a58554e",
  2261 => x"4f2c2041",
  2262 => x"454f4e2c",
  2263 => x"00000000",
  2264 => x"5a58444f",
  2265 => x"5320616e",
  2266 => x"64205a58",
  2267 => x"444f532b",
  2268 => x"20626f61",
  2269 => x"7264732e",
  2270 => x"00000000",
  2271 => x"4f726967",
  2272 => x"696e616c",
  2273 => x"20636f72",
  2274 => x"65206279",
  2275 => x"3a000000",
  2276 => x"202d2043",
  2277 => x"61727374",
  2278 => x"656e2045",
  2279 => x"6c746f6e",
  2280 => x"20536f72",
  2281 => x"656e7365",
  2282 => x"6e200000",
  2283 => x"506f7274",
  2284 => x"206d6164",
  2285 => x"65206279",
  2286 => x"3a000000",
  2287 => x"202d2041",
  2288 => x"7a65736d",
  2289 => x"626f6700",
  2290 => x"202d2041",
  2291 => x"766c6978",
  2292 => x"41000000",
  2293 => x"496e6974",
  2294 => x"69616c69",
  2295 => x"7a696e67",
  2296 => x"20534420",
  2297 => x"63617264",
  2298 => x"0a000000",
  2299 => x"5a583831",
  2300 => x"20202020",
  2301 => x"20202000",
  2302 => x"524f4d53",
  2303 => x"20202020",
  2304 => x"20202000",
  2305 => x"5a583858",
  2306 => x"20202020",
  2307 => x"524f4d00",
  2308 => x"4572726f",
  2309 => x"72204c6f",
  2310 => x"6164696e",
  2311 => x"6720524f",
  2312 => x"4d2e2e2e",
  2313 => x"0a000000",
  2314 => x"16200000",
  2315 => x"14200000",
  2316 => x"15200000",
  2317 => x"53442069",
  2318 => x"6e69742e",
  2319 => x"2e2e0a00",
  2320 => x"53442063",
  2321 => x"61726420",
  2322 => x"72657365",
  2323 => x"74206661",
  2324 => x"696c6564",
  2325 => x"210a0000",
  2326 => x"53444843",
  2327 => x"20657272",
  2328 => x"6f72210a",
  2329 => x"00000000",
  2330 => x"57726974",
  2331 => x"65206661",
  2332 => x"696c6564",
  2333 => x"0a000000",
  2334 => x"52656164",
  2335 => x"20666169",
  2336 => x"6c65640a",
  2337 => x"00000000",
  2338 => x"43617264",
  2339 => x"20696e69",
  2340 => x"74206661",
  2341 => x"696c6564",
  2342 => x"0a000000",
  2343 => x"46415431",
  2344 => x"36202020",
  2345 => x"00000000",
  2346 => x"46415433",
  2347 => x"32202020",
  2348 => x"00000000",
  2349 => x"4e6f2070",
  2350 => x"61727469",
  2351 => x"74696f6e",
  2352 => x"20736967",
  2353 => x"0a000000",
  2354 => x"42616420",
  2355 => x"70617274",
  2356 => x"0a000000",
  2357 => x"4261636b",
  2358 => x"00000000",
  2359 => x"00000002",
  2360 => x"00000002",
  2361 => x"00001ea4",
  2362 => x"0000036b",
  2363 => x"00000002",
  2364 => x"00001ec0",
  2365 => x"0000036b",
  2366 => x"00000003",
  2367 => x"000025cc",
  2368 => x"00000002",
  2369 => x"00000003",
  2370 => x"000025bc",
  2371 => x"00000004",
  2372 => x"00000001",
  2373 => x"00001edc",
  2374 => x"00000000",
  2375 => x"00000003",
  2376 => x"000025b0",
  2377 => x"00000003",
  2378 => x"00000001",
  2379 => x"00001ef0",
  2380 => x"00000001",
  2381 => x"00000003",
  2382 => x"000025a4",
  2383 => x"00000003",
  2384 => x"00000001",
  2385 => x"00001f10",
  2386 => x"00000002",
  2387 => x"00000001",
  2388 => x"00001f2c",
  2389 => x"00000003",
  2390 => x"00000001",
  2391 => x"00001f44",
  2392 => x"00000004",
  2393 => x"00000003",
  2394 => x"00002594",
  2395 => x"00000003",
  2396 => x"00000001",
  2397 => x"00001f5c",
  2398 => x"00000005",
  2399 => x"00000004",
  2400 => x"00001f78",
  2401 => x"00002968",
  2402 => x"00000000",
  2403 => x"00000000",
  2404 => x"00000000",
  2405 => x"00001f80",
  2406 => x"00001f9c",
  2407 => x"00001fb4",
  2408 => x"00001fc8",
  2409 => x"00001fdc",
  2410 => x"00001ff4",
  2411 => x"0000200c",
  2412 => x"00002024",
  2413 => x"00002038",
  2414 => x"0000204c",
  2415 => x"0000205c",
  2416 => x"0000206c",
  2417 => x"0000207c",
  2418 => x"0000208c",
  2419 => x"0000209c",
  2420 => x"000020b4",
  2421 => x"00000002",
  2422 => x"000020cc",
  2423 => x"0000036c",
  2424 => x"00000002",
  2425 => x"000020e8",
  2426 => x"0000036c",
  2427 => x"00000002",
  2428 => x"00002104",
  2429 => x"000003af",
  2430 => x"00000002",
  2431 => x"0000210c",
  2432 => x"00001e3f",
  2433 => x"00000002",
  2434 => x"00002120",
  2435 => x"00001e5f",
  2436 => x"00000002",
  2437 => x"00002134",
  2438 => x"0000037c",
  2439 => x"00000002",
  2440 => x"0000214c",
  2441 => x"0000038c",
  2442 => x"00000002",
  2443 => x"0000215c",
  2444 => x"00000919",
  2445 => x"00000000",
  2446 => x"00000000",
  2447 => x"00000000",
  2448 => x"00000004",
  2449 => x"00002164",
  2450 => x"00002640",
  2451 => x"00000004",
  2452 => x"00002178",
  2453 => x"00002968",
  2454 => x"00000000",
  2455 => x"00000000",
  2456 => x"00000000",
  2457 => x"00000004",
  2458 => x"0000217c",
  2459 => x"00002664",
  2460 => x"00000004",
  2461 => x"00002190",
  2462 => x"00002664",
  2463 => x"00000004",
  2464 => x"000021b0",
  2465 => x"00002664",
  2466 => x"00000004",
  2467 => x"000021cc",
  2468 => x"00002664",
  2469 => x"00000004",
  2470 => x"00002464",
  2471 => x"00002664",
  2472 => x"00000004",
  2473 => x"00001e98",
  2474 => x"00002968",
  2475 => x"00000000",
  2476 => x"00000000",
  2477 => x"00000000",
  2478 => x"00000002",
  2479 => x"00002204",
  2480 => x"0000036b",
  2481 => x"00000002",
  2482 => x"00001ec0",
  2483 => x"0000036b",
  2484 => x"00000002",
  2485 => x"00002220",
  2486 => x"0000036b",
  2487 => x"00000002",
  2488 => x"0000223c",
  2489 => x"0000036b",
  2490 => x"00000002",
  2491 => x"00002254",
  2492 => x"0000036b",
  2493 => x"00000002",
  2494 => x"00002270",
  2495 => x"0000036b",
  2496 => x"00000002",
  2497 => x"00002290",
  2498 => x"0000036b",
  2499 => x"00000002",
  2500 => x"000022b0",
  2501 => x"0000036b",
  2502 => x"00000002",
  2503 => x"000022cc",
  2504 => x"0000036b",
  2505 => x"00000002",
  2506 => x"000022ec",
  2507 => x"0000036b",
  2508 => x"00000002",
  2509 => x"00002304",
  2510 => x"0000036b",
  2511 => x"00000002",
  2512 => x"00002464",
  2513 => x"0000036b",
  2514 => x"00000004",
  2515 => x"00002178",
  2516 => x"00002968",
  2517 => x"00000000",
  2518 => x"00000000",
  2519 => x"00000000",
  2520 => x"00000002",
  2521 => x"00002324",
  2522 => x"0000036b",
  2523 => x"00000002",
  2524 => x"00001ec0",
  2525 => x"0000036b",
  2526 => x"00000002",
  2527 => x"00002340",
  2528 => x"0000036b",
  2529 => x"00000002",
  2530 => x"00002360",
  2531 => x"0000036b",
  2532 => x"00000002",
  2533 => x"00002464",
  2534 => x"0000036b",
  2535 => x"00000002",
  2536 => x"0000237c",
  2537 => x"0000036b",
  2538 => x"00000002",
  2539 => x"00002390",
  2540 => x"0000036b",
  2541 => x"00000002",
  2542 => x"00002464",
  2543 => x"0000036b",
  2544 => x"00000002",
  2545 => x"000023ac",
  2546 => x"0000036b",
  2547 => x"00000002",
  2548 => x"000023bc",
  2549 => x"0000036b",
  2550 => x"00000002",
  2551 => x"000023c8",
  2552 => x"0000036b",
  2553 => x"00000002",
  2554 => x"00002464",
  2555 => x"0000036b",
  2556 => x"00000004",
  2557 => x"00002178",
  2558 => x"00002968",
  2559 => x"00000000",
  2560 => x"00000000",
  2561 => x"00000000",
  2562 => x"00000000",
  2563 => x"00000000",
  2564 => x"00000000",
  2565 => x"00000000",
  2566 => x"00000000",
  2567 => x"00000000",
  2568 => x"00000000",
  2569 => x"00000000",
  2570 => x"00000000",
  2571 => x"00000000",
  2572 => x"00000000",
  2573 => x"00000000",
  2574 => x"00000000",
  2575 => x"00000000",
  2576 => x"00000000",
  2577 => x"00000000",
  2578 => x"00000000",
  2579 => x"00000000",
  2580 => x"00000006",
  2581 => x"00000043",
  2582 => x"00000042",
  2583 => x"0000003b",
  2584 => x"0000004b",
  2585 => x"0000007e",
  2586 => x"00000003",
  2587 => x"0000000b",
  2588 => x"00000083",
  2589 => x"00000023",
  2590 => x"0000007e",
  2591 => x"00000000",
  2592 => x"00000000",
  2593 => x"00000002",
  2594 => x"00002cf4",
  2595 => x"00001bf3",
  2596 => x"00000002",
  2597 => x"00002d12",
  2598 => x"00001bf3",
  2599 => x"00000002",
  2600 => x"00002d30",
  2601 => x"00001bf3",
  2602 => x"00000002",
  2603 => x"00002d4e",
  2604 => x"00001bf3",
  2605 => x"00000002",
  2606 => x"00002d6c",
  2607 => x"00001bf3",
  2608 => x"00000002",
  2609 => x"00002d8a",
  2610 => x"00001bf3",
  2611 => x"00000002",
  2612 => x"00002da8",
  2613 => x"00001bf3",
  2614 => x"00000002",
  2615 => x"00002dc6",
  2616 => x"00001bf3",
  2617 => x"00000002",
  2618 => x"00002de4",
  2619 => x"00001bf3",
  2620 => x"00000002",
  2621 => x"00002e02",
  2622 => x"00001bf3",
  2623 => x"00000002",
  2624 => x"00002e20",
  2625 => x"00001bf3",
  2626 => x"00000002",
  2627 => x"00002e3e",
  2628 => x"00001bf3",
  2629 => x"00000002",
  2630 => x"00002e5c",
  2631 => x"00001bf3",
  2632 => x"00000004",
  2633 => x"000024d4",
  2634 => x"00000000",
  2635 => x"00000000",
  2636 => x"00000000",
  2637 => x"00001da5",
  2638 => x"00000000",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memAWriteEnable = '1') and (from_zpu.memBWriteEnable = '1') and (from_zpu.memAAddr=from_zpu.memBAddr) and (from_zpu.memAWrite/=from_zpu.memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (from_zpu.memAWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memAWrite;
			to_zpu.memARead <= from_zpu.memAWrite;
		else
			to_zpu.memARead <= ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memBWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memBWrite;
			to_zpu.memBRead <= from_zpu.memBWrite;
		else
			to_zpu.memBRead <= ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;


end arch;

